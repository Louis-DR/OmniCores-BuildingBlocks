
`define INFINITE (1/0)

localparam bool true  = 1'b1;
localparam bool false = 1'b0;
