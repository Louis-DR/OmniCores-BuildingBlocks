// ╔═══════════════════════════════════════════════════════════════════════════╗
// ║ Project:     OmniCores-BuildingBlocks                                     ║
// ║ Author:      Louis Duret-Robert - louisduret@gmail.com                    ║
// ║ Website:     louis-dr.github.io                                           ║
// ║ License:     MIT License                                                  ║
// ║ File:        shifter_right.tb.sv                                          ║
// ╟───────────────────────────────────────────────────────────────────────────╢
// ║ This file is generated from the template shifter_right.tb.sv.j2 by J2GPP. ║
// ║ Do not edit it directly.                                                  ║
// ╟───────────────────────────────────────────────────────────────────────────╢
// ║ Description: Top-level testbench for the static right shifter.            ║
// ║                                                                           ║
// ╚═══════════════════════════════════════════════════════════════════════════╝



`timescale 1ns/1ns



module shifter_right_tb ();


logic start__shifter_right_tc__width_1__shift_0__pad_0;

logic start__shifter_right_tc__width_1__shift_1__pad_0;

logic start__shifter_right_tc__width_1__shift_0__pad_1;

logic start__shifter_right_tc__width_1__shift_1__pad_1;

logic start__shifter_right_tc__width_2__shift_0__pad_0;

logic start__shifter_right_tc__width_2__shift_1__pad_0;

logic start__shifter_right_tc__width_2__shift_2__pad_0;

logic start__shifter_right_tc__width_2__shift_3__pad_0;

logic start__shifter_right_tc__width_2__shift_0__pad_1;

logic start__shifter_right_tc__width_2__shift_1__pad_1;

logic start__shifter_right_tc__width_2__shift_2__pad_1;

logic start__shifter_right_tc__width_2__shift_3__pad_1;

logic start__shifter_right_tc__width_3__shift_0__pad_0;

logic start__shifter_right_tc__width_3__shift_1__pad_0;

logic start__shifter_right_tc__width_3__shift_2__pad_0;

logic start__shifter_right_tc__width_3__shift_3__pad_0;

logic start__shifter_right_tc__width_3__shift_4__pad_0;

logic start__shifter_right_tc__width_3__shift_5__pad_0;

logic start__shifter_right_tc__width_3__shift_0__pad_1;

logic start__shifter_right_tc__width_3__shift_1__pad_1;

logic start__shifter_right_tc__width_3__shift_2__pad_1;

logic start__shifter_right_tc__width_3__shift_3__pad_1;

logic start__shifter_right_tc__width_3__shift_4__pad_1;

logic start__shifter_right_tc__width_3__shift_5__pad_1;

logic start__shifter_right_tc__width_4__shift_0__pad_0;

logic start__shifter_right_tc__width_4__shift_1__pad_0;

logic start__shifter_right_tc__width_4__shift_2__pad_0;

logic start__shifter_right_tc__width_4__shift_3__pad_0;

logic start__shifter_right_tc__width_4__shift_4__pad_0;

logic start__shifter_right_tc__width_4__shift_5__pad_0;

logic start__shifter_right_tc__width_4__shift_6__pad_0;

logic start__shifter_right_tc__width_4__shift_7__pad_0;

logic start__shifter_right_tc__width_4__shift_0__pad_1;

logic start__shifter_right_tc__width_4__shift_1__pad_1;

logic start__shifter_right_tc__width_4__shift_2__pad_1;

logic start__shifter_right_tc__width_4__shift_3__pad_1;

logic start__shifter_right_tc__width_4__shift_4__pad_1;

logic start__shifter_right_tc__width_4__shift_5__pad_1;

logic start__shifter_right_tc__width_4__shift_6__pad_1;

logic start__shifter_right_tc__width_4__shift_7__pad_1;

logic start__shifter_right_tc__width_5__shift_0__pad_0;

logic start__shifter_right_tc__width_5__shift_1__pad_0;

logic start__shifter_right_tc__width_5__shift_2__pad_0;

logic start__shifter_right_tc__width_5__shift_3__pad_0;

logic start__shifter_right_tc__width_5__shift_4__pad_0;

logic start__shifter_right_tc__width_5__shift_5__pad_0;

logic start__shifter_right_tc__width_5__shift_6__pad_0;

logic start__shifter_right_tc__width_5__shift_7__pad_0;

logic start__shifter_right_tc__width_5__shift_8__pad_0;

logic start__shifter_right_tc__width_5__shift_9__pad_0;

logic start__shifter_right_tc__width_5__shift_0__pad_1;

logic start__shifter_right_tc__width_5__shift_1__pad_1;

logic start__shifter_right_tc__width_5__shift_2__pad_1;

logic start__shifter_right_tc__width_5__shift_3__pad_1;

logic start__shifter_right_tc__width_5__shift_4__pad_1;

logic start__shifter_right_tc__width_5__shift_5__pad_1;

logic start__shifter_right_tc__width_5__shift_6__pad_1;

logic start__shifter_right_tc__width_5__shift_7__pad_1;

logic start__shifter_right_tc__width_5__shift_8__pad_1;

logic start__shifter_right_tc__width_5__shift_9__pad_1;

logic start__shifter_right_tc__width_6__shift_0__pad_0;

logic start__shifter_right_tc__width_6__shift_1__pad_0;

logic start__shifter_right_tc__width_6__shift_2__pad_0;

logic start__shifter_right_tc__width_6__shift_3__pad_0;

logic start__shifter_right_tc__width_6__shift_4__pad_0;

logic start__shifter_right_tc__width_6__shift_5__pad_0;

logic start__shifter_right_tc__width_6__shift_6__pad_0;

logic start__shifter_right_tc__width_6__shift_7__pad_0;

logic start__shifter_right_tc__width_6__shift_8__pad_0;

logic start__shifter_right_tc__width_6__shift_9__pad_0;

logic start__shifter_right_tc__width_6__shift_10__pad_0;

logic start__shifter_right_tc__width_6__shift_11__pad_0;

logic start__shifter_right_tc__width_6__shift_0__pad_1;

logic start__shifter_right_tc__width_6__shift_1__pad_1;

logic start__shifter_right_tc__width_6__shift_2__pad_1;

logic start__shifter_right_tc__width_6__shift_3__pad_1;

logic start__shifter_right_tc__width_6__shift_4__pad_1;

logic start__shifter_right_tc__width_6__shift_5__pad_1;

logic start__shifter_right_tc__width_6__shift_6__pad_1;

logic start__shifter_right_tc__width_6__shift_7__pad_1;

logic start__shifter_right_tc__width_6__shift_8__pad_1;

logic start__shifter_right_tc__width_6__shift_9__pad_1;

logic start__shifter_right_tc__width_6__shift_10__pad_1;

logic start__shifter_right_tc__width_6__shift_11__pad_1;

logic start__shifter_right_tc__width_7__shift_0__pad_0;

logic start__shifter_right_tc__width_7__shift_1__pad_0;

logic start__shifter_right_tc__width_7__shift_2__pad_0;

logic start__shifter_right_tc__width_7__shift_3__pad_0;

logic start__shifter_right_tc__width_7__shift_4__pad_0;

logic start__shifter_right_tc__width_7__shift_5__pad_0;

logic start__shifter_right_tc__width_7__shift_6__pad_0;

logic start__shifter_right_tc__width_7__shift_7__pad_0;

logic start__shifter_right_tc__width_7__shift_8__pad_0;

logic start__shifter_right_tc__width_7__shift_9__pad_0;

logic start__shifter_right_tc__width_7__shift_10__pad_0;

logic start__shifter_right_tc__width_7__shift_11__pad_0;

logic start__shifter_right_tc__width_7__shift_12__pad_0;

logic start__shifter_right_tc__width_7__shift_13__pad_0;

logic start__shifter_right_tc__width_7__shift_0__pad_1;

logic start__shifter_right_tc__width_7__shift_1__pad_1;

logic start__shifter_right_tc__width_7__shift_2__pad_1;

logic start__shifter_right_tc__width_7__shift_3__pad_1;

logic start__shifter_right_tc__width_7__shift_4__pad_1;

logic start__shifter_right_tc__width_7__shift_5__pad_1;

logic start__shifter_right_tc__width_7__shift_6__pad_1;

logic start__shifter_right_tc__width_7__shift_7__pad_1;

logic start__shifter_right_tc__width_7__shift_8__pad_1;

logic start__shifter_right_tc__width_7__shift_9__pad_1;

logic start__shifter_right_tc__width_7__shift_10__pad_1;

logic start__shifter_right_tc__width_7__shift_11__pad_1;

logic start__shifter_right_tc__width_7__shift_12__pad_1;

logic start__shifter_right_tc__width_7__shift_13__pad_1;

logic start__shifter_right_tc__width_8__shift_0__pad_0;

logic start__shifter_right_tc__width_8__shift_1__pad_0;

logic start__shifter_right_tc__width_8__shift_2__pad_0;

logic start__shifter_right_tc__width_8__shift_3__pad_0;

logic start__shifter_right_tc__width_8__shift_4__pad_0;

logic start__shifter_right_tc__width_8__shift_5__pad_0;

logic start__shifter_right_tc__width_8__shift_6__pad_0;

logic start__shifter_right_tc__width_8__shift_7__pad_0;

logic start__shifter_right_tc__width_8__shift_8__pad_0;

logic start__shifter_right_tc__width_8__shift_9__pad_0;

logic start__shifter_right_tc__width_8__shift_10__pad_0;

logic start__shifter_right_tc__width_8__shift_11__pad_0;

logic start__shifter_right_tc__width_8__shift_12__pad_0;

logic start__shifter_right_tc__width_8__shift_13__pad_0;

logic start__shifter_right_tc__width_8__shift_14__pad_0;

logic start__shifter_right_tc__width_8__shift_15__pad_0;

logic start__shifter_right_tc__width_8__shift_0__pad_1;

logic start__shifter_right_tc__width_8__shift_1__pad_1;

logic start__shifter_right_tc__width_8__shift_2__pad_1;

logic start__shifter_right_tc__width_8__shift_3__pad_1;

logic start__shifter_right_tc__width_8__shift_4__pad_1;

logic start__shifter_right_tc__width_8__shift_5__pad_1;

logic start__shifter_right_tc__width_8__shift_6__pad_1;

logic start__shifter_right_tc__width_8__shift_7__pad_1;

logic start__shifter_right_tc__width_8__shift_8__pad_1;

logic start__shifter_right_tc__width_8__shift_9__pad_1;

logic start__shifter_right_tc__width_8__shift_10__pad_1;

logic start__shifter_right_tc__width_8__shift_11__pad_1;

logic start__shifter_right_tc__width_8__shift_12__pad_1;

logic start__shifter_right_tc__width_8__shift_13__pad_1;

logic start__shifter_right_tc__width_8__shift_14__pad_1;

logic start__shifter_right_tc__width_8__shift_15__pad_1;

logic start__shifter_right_tc__width_9__shift_0__pad_0;

logic start__shifter_right_tc__width_9__shift_1__pad_0;

logic start__shifter_right_tc__width_9__shift_2__pad_0;

logic start__shifter_right_tc__width_9__shift_3__pad_0;

logic start__shifter_right_tc__width_9__shift_4__pad_0;

logic start__shifter_right_tc__width_9__shift_5__pad_0;

logic start__shifter_right_tc__width_9__shift_6__pad_0;

logic start__shifter_right_tc__width_9__shift_7__pad_0;

logic start__shifter_right_tc__width_9__shift_8__pad_0;

logic start__shifter_right_tc__width_9__shift_9__pad_0;

logic start__shifter_right_tc__width_9__shift_10__pad_0;

logic start__shifter_right_tc__width_9__shift_11__pad_0;

logic start__shifter_right_tc__width_9__shift_12__pad_0;

logic start__shifter_right_tc__width_9__shift_13__pad_0;

logic start__shifter_right_tc__width_9__shift_14__pad_0;

logic start__shifter_right_tc__width_9__shift_15__pad_0;

logic start__shifter_right_tc__width_9__shift_16__pad_0;

logic start__shifter_right_tc__width_9__shift_17__pad_0;

logic start__shifter_right_tc__width_9__shift_0__pad_1;

logic start__shifter_right_tc__width_9__shift_1__pad_1;

logic start__shifter_right_tc__width_9__shift_2__pad_1;

logic start__shifter_right_tc__width_9__shift_3__pad_1;

logic start__shifter_right_tc__width_9__shift_4__pad_1;

logic start__shifter_right_tc__width_9__shift_5__pad_1;

logic start__shifter_right_tc__width_9__shift_6__pad_1;

logic start__shifter_right_tc__width_9__shift_7__pad_1;

logic start__shifter_right_tc__width_9__shift_8__pad_1;

logic start__shifter_right_tc__width_9__shift_9__pad_1;

logic start__shifter_right_tc__width_9__shift_10__pad_1;

logic start__shifter_right_tc__width_9__shift_11__pad_1;

logic start__shifter_right_tc__width_9__shift_12__pad_1;

logic start__shifter_right_tc__width_9__shift_13__pad_1;

logic start__shifter_right_tc__width_9__shift_14__pad_1;

logic start__shifter_right_tc__width_9__shift_15__pad_1;

logic start__shifter_right_tc__width_9__shift_16__pad_1;

logic start__shifter_right_tc__width_9__shift_17__pad_1;

logic start__shifter_right_tc__width_10__shift_0__pad_0;

logic start__shifter_right_tc__width_10__shift_1__pad_0;

logic start__shifter_right_tc__width_10__shift_2__pad_0;

logic start__shifter_right_tc__width_10__shift_3__pad_0;

logic start__shifter_right_tc__width_10__shift_4__pad_0;

logic start__shifter_right_tc__width_10__shift_5__pad_0;

logic start__shifter_right_tc__width_10__shift_6__pad_0;

logic start__shifter_right_tc__width_10__shift_7__pad_0;

logic start__shifter_right_tc__width_10__shift_8__pad_0;

logic start__shifter_right_tc__width_10__shift_9__pad_0;

logic start__shifter_right_tc__width_10__shift_10__pad_0;

logic start__shifter_right_tc__width_10__shift_11__pad_0;

logic start__shifter_right_tc__width_10__shift_12__pad_0;

logic start__shifter_right_tc__width_10__shift_13__pad_0;

logic start__shifter_right_tc__width_10__shift_14__pad_0;

logic start__shifter_right_tc__width_10__shift_15__pad_0;

logic start__shifter_right_tc__width_10__shift_16__pad_0;

logic start__shifter_right_tc__width_10__shift_17__pad_0;

logic start__shifter_right_tc__width_10__shift_18__pad_0;

logic start__shifter_right_tc__width_10__shift_19__pad_0;

logic start__shifter_right_tc__width_10__shift_0__pad_1;

logic start__shifter_right_tc__width_10__shift_1__pad_1;

logic start__shifter_right_tc__width_10__shift_2__pad_1;

logic start__shifter_right_tc__width_10__shift_3__pad_1;

logic start__shifter_right_tc__width_10__shift_4__pad_1;

logic start__shifter_right_tc__width_10__shift_5__pad_1;

logic start__shifter_right_tc__width_10__shift_6__pad_1;

logic start__shifter_right_tc__width_10__shift_7__pad_1;

logic start__shifter_right_tc__width_10__shift_8__pad_1;

logic start__shifter_right_tc__width_10__shift_9__pad_1;

logic start__shifter_right_tc__width_10__shift_10__pad_1;

logic start__shifter_right_tc__width_10__shift_11__pad_1;

logic start__shifter_right_tc__width_10__shift_12__pad_1;

logic start__shifter_right_tc__width_10__shift_13__pad_1;

logic start__shifter_right_tc__width_10__shift_14__pad_1;

logic start__shifter_right_tc__width_10__shift_15__pad_1;

logic start__shifter_right_tc__width_10__shift_16__pad_1;

logic start__shifter_right_tc__width_10__shift_17__pad_1;

logic start__shifter_right_tc__width_10__shift_18__pad_1;

logic start__shifter_right_tc__width_10__shift_19__pad_1;

logic start__shifter_right_tc__width_11__shift_0__pad_0;

logic start__shifter_right_tc__width_11__shift_1__pad_0;

logic start__shifter_right_tc__width_11__shift_2__pad_0;

logic start__shifter_right_tc__width_11__shift_3__pad_0;

logic start__shifter_right_tc__width_11__shift_4__pad_0;

logic start__shifter_right_tc__width_11__shift_5__pad_0;

logic start__shifter_right_tc__width_11__shift_6__pad_0;

logic start__shifter_right_tc__width_11__shift_7__pad_0;

logic start__shifter_right_tc__width_11__shift_8__pad_0;

logic start__shifter_right_tc__width_11__shift_9__pad_0;

logic start__shifter_right_tc__width_11__shift_10__pad_0;

logic start__shifter_right_tc__width_11__shift_11__pad_0;

logic start__shifter_right_tc__width_11__shift_12__pad_0;

logic start__shifter_right_tc__width_11__shift_13__pad_0;

logic start__shifter_right_tc__width_11__shift_14__pad_0;

logic start__shifter_right_tc__width_11__shift_15__pad_0;

logic start__shifter_right_tc__width_11__shift_16__pad_0;

logic start__shifter_right_tc__width_11__shift_17__pad_0;

logic start__shifter_right_tc__width_11__shift_18__pad_0;

logic start__shifter_right_tc__width_11__shift_19__pad_0;

logic start__shifter_right_tc__width_11__shift_20__pad_0;

logic start__shifter_right_tc__width_11__shift_21__pad_0;

logic start__shifter_right_tc__width_11__shift_0__pad_1;

logic start__shifter_right_tc__width_11__shift_1__pad_1;

logic start__shifter_right_tc__width_11__shift_2__pad_1;

logic start__shifter_right_tc__width_11__shift_3__pad_1;

logic start__shifter_right_tc__width_11__shift_4__pad_1;

logic start__shifter_right_tc__width_11__shift_5__pad_1;

logic start__shifter_right_tc__width_11__shift_6__pad_1;

logic start__shifter_right_tc__width_11__shift_7__pad_1;

logic start__shifter_right_tc__width_11__shift_8__pad_1;

logic start__shifter_right_tc__width_11__shift_9__pad_1;

logic start__shifter_right_tc__width_11__shift_10__pad_1;

logic start__shifter_right_tc__width_11__shift_11__pad_1;

logic start__shifter_right_tc__width_11__shift_12__pad_1;

logic start__shifter_right_tc__width_11__shift_13__pad_1;

logic start__shifter_right_tc__width_11__shift_14__pad_1;

logic start__shifter_right_tc__width_11__shift_15__pad_1;

logic start__shifter_right_tc__width_11__shift_16__pad_1;

logic start__shifter_right_tc__width_11__shift_17__pad_1;

logic start__shifter_right_tc__width_11__shift_18__pad_1;

logic start__shifter_right_tc__width_11__shift_19__pad_1;

logic start__shifter_right_tc__width_11__shift_20__pad_1;

logic start__shifter_right_tc__width_11__shift_21__pad_1;

logic start__shifter_right_tc__width_12__shift_0__pad_0;

logic start__shifter_right_tc__width_12__shift_1__pad_0;

logic start__shifter_right_tc__width_12__shift_2__pad_0;

logic start__shifter_right_tc__width_12__shift_3__pad_0;

logic start__shifter_right_tc__width_12__shift_4__pad_0;

logic start__shifter_right_tc__width_12__shift_5__pad_0;

logic start__shifter_right_tc__width_12__shift_6__pad_0;

logic start__shifter_right_tc__width_12__shift_7__pad_0;

logic start__shifter_right_tc__width_12__shift_8__pad_0;

logic start__shifter_right_tc__width_12__shift_9__pad_0;

logic start__shifter_right_tc__width_12__shift_10__pad_0;

logic start__shifter_right_tc__width_12__shift_11__pad_0;

logic start__shifter_right_tc__width_12__shift_12__pad_0;

logic start__shifter_right_tc__width_12__shift_13__pad_0;

logic start__shifter_right_tc__width_12__shift_14__pad_0;

logic start__shifter_right_tc__width_12__shift_15__pad_0;

logic start__shifter_right_tc__width_12__shift_16__pad_0;

logic start__shifter_right_tc__width_12__shift_17__pad_0;

logic start__shifter_right_tc__width_12__shift_18__pad_0;

logic start__shifter_right_tc__width_12__shift_19__pad_0;

logic start__shifter_right_tc__width_12__shift_20__pad_0;

logic start__shifter_right_tc__width_12__shift_21__pad_0;

logic start__shifter_right_tc__width_12__shift_22__pad_0;

logic start__shifter_right_tc__width_12__shift_23__pad_0;

logic start__shifter_right_tc__width_12__shift_0__pad_1;

logic start__shifter_right_tc__width_12__shift_1__pad_1;

logic start__shifter_right_tc__width_12__shift_2__pad_1;

logic start__shifter_right_tc__width_12__shift_3__pad_1;

logic start__shifter_right_tc__width_12__shift_4__pad_1;

logic start__shifter_right_tc__width_12__shift_5__pad_1;

logic start__shifter_right_tc__width_12__shift_6__pad_1;

logic start__shifter_right_tc__width_12__shift_7__pad_1;

logic start__shifter_right_tc__width_12__shift_8__pad_1;

logic start__shifter_right_tc__width_12__shift_9__pad_1;

logic start__shifter_right_tc__width_12__shift_10__pad_1;

logic start__shifter_right_tc__width_12__shift_11__pad_1;

logic start__shifter_right_tc__width_12__shift_12__pad_1;

logic start__shifter_right_tc__width_12__shift_13__pad_1;

logic start__shifter_right_tc__width_12__shift_14__pad_1;

logic start__shifter_right_tc__width_12__shift_15__pad_1;

logic start__shifter_right_tc__width_12__shift_16__pad_1;

logic start__shifter_right_tc__width_12__shift_17__pad_1;

logic start__shifter_right_tc__width_12__shift_18__pad_1;

logic start__shifter_right_tc__width_12__shift_19__pad_1;

logic start__shifter_right_tc__width_12__shift_20__pad_1;

logic start__shifter_right_tc__width_12__shift_21__pad_1;

logic start__shifter_right_tc__width_12__shift_22__pad_1;

logic start__shifter_right_tc__width_12__shift_23__pad_1;

logic start__shifter_right_tc__width_16__shift_0__pad_0;

logic start__shifter_right_tc__width_16__shift_1__pad_0;

logic start__shifter_right_tc__width_16__shift_2__pad_0;

logic start__shifter_right_tc__width_16__shift_3__pad_0;

logic start__shifter_right_tc__width_16__shift_4__pad_0;

logic start__shifter_right_tc__width_16__shift_5__pad_0;

logic start__shifter_right_tc__width_16__shift_6__pad_0;

logic start__shifter_right_tc__width_16__shift_7__pad_0;

logic start__shifter_right_tc__width_16__shift_8__pad_0;

logic start__shifter_right_tc__width_16__shift_15__pad_0;

logic start__shifter_right_tc__width_16__shift_16__pad_0;

logic start__shifter_right_tc__width_16__shift_17__pad_0;

logic start__shifter_right_tc__width_16__shift_24__pad_0;

logic start__shifter_right_tc__width_16__shift_31__pad_0;

logic start__shifter_right_tc__width_16__shift_32__pad_0;

logic start__shifter_right_tc__width_16__shift_0__pad_1;

logic start__shifter_right_tc__width_16__shift_1__pad_1;

logic start__shifter_right_tc__width_16__shift_2__pad_1;

logic start__shifter_right_tc__width_16__shift_3__pad_1;

logic start__shifter_right_tc__width_16__shift_4__pad_1;

logic start__shifter_right_tc__width_16__shift_5__pad_1;

logic start__shifter_right_tc__width_16__shift_6__pad_1;

logic start__shifter_right_tc__width_16__shift_7__pad_1;

logic start__shifter_right_tc__width_16__shift_8__pad_1;

logic start__shifter_right_tc__width_16__shift_15__pad_1;

logic start__shifter_right_tc__width_16__shift_16__pad_1;

logic start__shifter_right_tc__width_16__shift_17__pad_1;

logic start__shifter_right_tc__width_16__shift_24__pad_1;

logic start__shifter_right_tc__width_16__shift_31__pad_1;

logic start__shifter_right_tc__width_16__shift_32__pad_1;

logic start__shifter_right_tc__width_24__shift_0__pad_0;

logic start__shifter_right_tc__width_24__shift_1__pad_0;

logic start__shifter_right_tc__width_24__shift_2__pad_0;

logic start__shifter_right_tc__width_24__shift_3__pad_0;

logic start__shifter_right_tc__width_24__shift_4__pad_0;

logic start__shifter_right_tc__width_24__shift_5__pad_0;

logic start__shifter_right_tc__width_24__shift_6__pad_0;

logic start__shifter_right_tc__width_24__shift_7__pad_0;

logic start__shifter_right_tc__width_24__shift_12__pad_0;

logic start__shifter_right_tc__width_24__shift_23__pad_0;

logic start__shifter_right_tc__width_24__shift_24__pad_0;

logic start__shifter_right_tc__width_24__shift_25__pad_0;

logic start__shifter_right_tc__width_24__shift_36__pad_0;

logic start__shifter_right_tc__width_24__shift_47__pad_0;

logic start__shifter_right_tc__width_24__shift_48__pad_0;

logic start__shifter_right_tc__width_24__shift_0__pad_1;

logic start__shifter_right_tc__width_24__shift_1__pad_1;

logic start__shifter_right_tc__width_24__shift_2__pad_1;

logic start__shifter_right_tc__width_24__shift_3__pad_1;

logic start__shifter_right_tc__width_24__shift_4__pad_1;

logic start__shifter_right_tc__width_24__shift_5__pad_1;

logic start__shifter_right_tc__width_24__shift_6__pad_1;

logic start__shifter_right_tc__width_24__shift_7__pad_1;

logic start__shifter_right_tc__width_24__shift_12__pad_1;

logic start__shifter_right_tc__width_24__shift_23__pad_1;

logic start__shifter_right_tc__width_24__shift_24__pad_1;

logic start__shifter_right_tc__width_24__shift_25__pad_1;

logic start__shifter_right_tc__width_24__shift_36__pad_1;

logic start__shifter_right_tc__width_24__shift_47__pad_1;

logic start__shifter_right_tc__width_24__shift_48__pad_1;

logic start__shifter_right_tc__width_32__shift_0__pad_0;

logic start__shifter_right_tc__width_32__shift_1__pad_0;

logic start__shifter_right_tc__width_32__shift_2__pad_0;

logic start__shifter_right_tc__width_32__shift_3__pad_0;

logic start__shifter_right_tc__width_32__shift_4__pad_0;

logic start__shifter_right_tc__width_32__shift_5__pad_0;

logic start__shifter_right_tc__width_32__shift_6__pad_0;

logic start__shifter_right_tc__width_32__shift_7__pad_0;

logic start__shifter_right_tc__width_32__shift_16__pad_0;

logic start__shifter_right_tc__width_32__shift_31__pad_0;

logic start__shifter_right_tc__width_32__shift_32__pad_0;

logic start__shifter_right_tc__width_32__shift_33__pad_0;

logic start__shifter_right_tc__width_32__shift_48__pad_0;

logic start__shifter_right_tc__width_32__shift_63__pad_0;

logic start__shifter_right_tc__width_32__shift_64__pad_0;

logic start__shifter_right_tc__width_32__shift_0__pad_1;

logic start__shifter_right_tc__width_32__shift_1__pad_1;

logic start__shifter_right_tc__width_32__shift_2__pad_1;

logic start__shifter_right_tc__width_32__shift_3__pad_1;

logic start__shifter_right_tc__width_32__shift_4__pad_1;

logic start__shifter_right_tc__width_32__shift_5__pad_1;

logic start__shifter_right_tc__width_32__shift_6__pad_1;

logic start__shifter_right_tc__width_32__shift_7__pad_1;

logic start__shifter_right_tc__width_32__shift_16__pad_1;

logic start__shifter_right_tc__width_32__shift_31__pad_1;

logic start__shifter_right_tc__width_32__shift_32__pad_1;

logic start__shifter_right_tc__width_32__shift_33__pad_1;

logic start__shifter_right_tc__width_32__shift_48__pad_1;

logic start__shifter_right_tc__width_32__shift_63__pad_1;

logic start__shifter_right_tc__width_32__shift_64__pad_1;

logic start__shifter_right_tc__width_48__shift_0__pad_0;

logic start__shifter_right_tc__width_48__shift_1__pad_0;

logic start__shifter_right_tc__width_48__shift_2__pad_0;

logic start__shifter_right_tc__width_48__shift_3__pad_0;

logic start__shifter_right_tc__width_48__shift_4__pad_0;

logic start__shifter_right_tc__width_48__shift_5__pad_0;

logic start__shifter_right_tc__width_48__shift_6__pad_0;

logic start__shifter_right_tc__width_48__shift_7__pad_0;

logic start__shifter_right_tc__width_48__shift_24__pad_0;

logic start__shifter_right_tc__width_48__shift_47__pad_0;

logic start__shifter_right_tc__width_48__shift_48__pad_0;

logic start__shifter_right_tc__width_48__shift_49__pad_0;

logic start__shifter_right_tc__width_48__shift_72__pad_0;

logic start__shifter_right_tc__width_48__shift_95__pad_0;

logic start__shifter_right_tc__width_48__shift_96__pad_0;

logic start__shifter_right_tc__width_48__shift_0__pad_1;

logic start__shifter_right_tc__width_48__shift_1__pad_1;

logic start__shifter_right_tc__width_48__shift_2__pad_1;

logic start__shifter_right_tc__width_48__shift_3__pad_1;

logic start__shifter_right_tc__width_48__shift_4__pad_1;

logic start__shifter_right_tc__width_48__shift_5__pad_1;

logic start__shifter_right_tc__width_48__shift_6__pad_1;

logic start__shifter_right_tc__width_48__shift_7__pad_1;

logic start__shifter_right_tc__width_48__shift_24__pad_1;

logic start__shifter_right_tc__width_48__shift_47__pad_1;

logic start__shifter_right_tc__width_48__shift_48__pad_1;

logic start__shifter_right_tc__width_48__shift_49__pad_1;

logic start__shifter_right_tc__width_48__shift_72__pad_1;

logic start__shifter_right_tc__width_48__shift_95__pad_1;

logic start__shifter_right_tc__width_48__shift_96__pad_1;

logic start__shifter_right_tc__width_64__shift_0__pad_0;

logic start__shifter_right_tc__width_64__shift_1__pad_0;

logic start__shifter_right_tc__width_64__shift_2__pad_0;

logic start__shifter_right_tc__width_64__shift_3__pad_0;

logic start__shifter_right_tc__width_64__shift_4__pad_0;

logic start__shifter_right_tc__width_64__shift_5__pad_0;

logic start__shifter_right_tc__width_64__shift_6__pad_0;

logic start__shifter_right_tc__width_64__shift_7__pad_0;

logic start__shifter_right_tc__width_64__shift_32__pad_0;

logic start__shifter_right_tc__width_64__shift_63__pad_0;

logic start__shifter_right_tc__width_64__shift_64__pad_0;

logic start__shifter_right_tc__width_64__shift_65__pad_0;

logic start__shifter_right_tc__width_64__shift_96__pad_0;

logic start__shifter_right_tc__width_64__shift_127__pad_0;

logic start__shifter_right_tc__width_64__shift_128__pad_0;

logic start__shifter_right_tc__width_64__shift_0__pad_1;

logic start__shifter_right_tc__width_64__shift_1__pad_1;

logic start__shifter_right_tc__width_64__shift_2__pad_1;

logic start__shifter_right_tc__width_64__shift_3__pad_1;

logic start__shifter_right_tc__width_64__shift_4__pad_1;

logic start__shifter_right_tc__width_64__shift_5__pad_1;

logic start__shifter_right_tc__width_64__shift_6__pad_1;

logic start__shifter_right_tc__width_64__shift_7__pad_1;

logic start__shifter_right_tc__width_64__shift_32__pad_1;

logic start__shifter_right_tc__width_64__shift_63__pad_1;

logic start__shifter_right_tc__width_64__shift_64__pad_1;

logic start__shifter_right_tc__width_64__shift_65__pad_1;

logic start__shifter_right_tc__width_64__shift_96__pad_1;

logic start__shifter_right_tc__width_64__shift_127__pad_1;

logic start__shifter_right_tc__width_64__shift_128__pad_1;

logic start__shifter_right_tc__width_128__shift_0__pad_0;

logic start__shifter_right_tc__width_128__shift_1__pad_0;

logic start__shifter_right_tc__width_128__shift_2__pad_0;

logic start__shifter_right_tc__width_128__shift_3__pad_0;

logic start__shifter_right_tc__width_128__shift_4__pad_0;

logic start__shifter_right_tc__width_128__shift_5__pad_0;

logic start__shifter_right_tc__width_128__shift_6__pad_0;

logic start__shifter_right_tc__width_128__shift_7__pad_0;

logic start__shifter_right_tc__width_128__shift_64__pad_0;

logic start__shifter_right_tc__width_128__shift_127__pad_0;

logic start__shifter_right_tc__width_128__shift_128__pad_0;

logic start__shifter_right_tc__width_128__shift_129__pad_0;

logic start__shifter_right_tc__width_128__shift_192__pad_0;

logic start__shifter_right_tc__width_128__shift_255__pad_0;

logic start__shifter_right_tc__width_128__shift_256__pad_0;

logic start__shifter_right_tc__width_128__shift_0__pad_1;

logic start__shifter_right_tc__width_128__shift_1__pad_1;

logic start__shifter_right_tc__width_128__shift_2__pad_1;

logic start__shifter_right_tc__width_128__shift_3__pad_1;

logic start__shifter_right_tc__width_128__shift_4__pad_1;

logic start__shifter_right_tc__width_128__shift_5__pad_1;

logic start__shifter_right_tc__width_128__shift_6__pad_1;

logic start__shifter_right_tc__width_128__shift_7__pad_1;

logic start__shifter_right_tc__width_128__shift_64__pad_1;

logic start__shifter_right_tc__width_128__shift_127__pad_1;

logic start__shifter_right_tc__width_128__shift_128__pad_1;

logic start__shifter_right_tc__width_128__shift_129__pad_1;

logic start__shifter_right_tc__width_128__shift_192__pad_1;

logic start__shifter_right_tc__width_128__shift_255__pad_1;

logic start__shifter_right_tc__width_128__shift_256__pad_1;

logic start__shifter_right_tc__width_256__shift_0__pad_0;

logic start__shifter_right_tc__width_256__shift_1__pad_0;

logic start__shifter_right_tc__width_256__shift_2__pad_0;

logic start__shifter_right_tc__width_256__shift_3__pad_0;

logic start__shifter_right_tc__width_256__shift_4__pad_0;

logic start__shifter_right_tc__width_256__shift_5__pad_0;

logic start__shifter_right_tc__width_256__shift_6__pad_0;

logic start__shifter_right_tc__width_256__shift_7__pad_0;

logic start__shifter_right_tc__width_256__shift_128__pad_0;

logic start__shifter_right_tc__width_256__shift_255__pad_0;

logic start__shifter_right_tc__width_256__shift_256__pad_0;

logic start__shifter_right_tc__width_256__shift_257__pad_0;

logic start__shifter_right_tc__width_256__shift_384__pad_0;

logic start__shifter_right_tc__width_256__shift_511__pad_0;

logic start__shifter_right_tc__width_256__shift_512__pad_0;

logic start__shifter_right_tc__width_256__shift_0__pad_1;

logic start__shifter_right_tc__width_256__shift_1__pad_1;

logic start__shifter_right_tc__width_256__shift_2__pad_1;

logic start__shifter_right_tc__width_256__shift_3__pad_1;

logic start__shifter_right_tc__width_256__shift_4__pad_1;

logic start__shifter_right_tc__width_256__shift_5__pad_1;

logic start__shifter_right_tc__width_256__shift_6__pad_1;

logic start__shifter_right_tc__width_256__shift_7__pad_1;

logic start__shifter_right_tc__width_256__shift_128__pad_1;

logic start__shifter_right_tc__width_256__shift_255__pad_1;

logic start__shifter_right_tc__width_256__shift_256__pad_1;

logic start__shifter_right_tc__width_256__shift_257__pad_1;

logic start__shifter_right_tc__width_256__shift_384__pad_1;

logic start__shifter_right_tc__width_256__shift_511__pad_1;

logic start__shifter_right_tc__width_256__shift_512__pad_1;

logic start__shifter_right_tc__width_512__shift_0__pad_0;

logic start__shifter_right_tc__width_512__shift_1__pad_0;

logic start__shifter_right_tc__width_512__shift_2__pad_0;

logic start__shifter_right_tc__width_512__shift_3__pad_0;

logic start__shifter_right_tc__width_512__shift_4__pad_0;

logic start__shifter_right_tc__width_512__shift_5__pad_0;

logic start__shifter_right_tc__width_512__shift_6__pad_0;

logic start__shifter_right_tc__width_512__shift_7__pad_0;

logic start__shifter_right_tc__width_512__shift_256__pad_0;

logic start__shifter_right_tc__width_512__shift_511__pad_0;

logic start__shifter_right_tc__width_512__shift_512__pad_0;

logic start__shifter_right_tc__width_512__shift_513__pad_0;

logic start__shifter_right_tc__width_512__shift_768__pad_0;

logic start__shifter_right_tc__width_512__shift_1023__pad_0;

logic start__shifter_right_tc__width_512__shift_1024__pad_0;

logic start__shifter_right_tc__width_512__shift_0__pad_1;

logic start__shifter_right_tc__width_512__shift_1__pad_1;

logic start__shifter_right_tc__width_512__shift_2__pad_1;

logic start__shifter_right_tc__width_512__shift_3__pad_1;

logic start__shifter_right_tc__width_512__shift_4__pad_1;

logic start__shifter_right_tc__width_512__shift_5__pad_1;

logic start__shifter_right_tc__width_512__shift_6__pad_1;

logic start__shifter_right_tc__width_512__shift_7__pad_1;

logic start__shifter_right_tc__width_512__shift_256__pad_1;

logic start__shifter_right_tc__width_512__shift_511__pad_1;

logic start__shifter_right_tc__width_512__shift_512__pad_1;

logic start__shifter_right_tc__width_512__shift_513__pad_1;

logic start__shifter_right_tc__width_512__shift_768__pad_1;

logic start__shifter_right_tc__width_512__shift_1023__pad_1;

logic start__shifter_right_tc__width_512__shift_1024__pad_1;

logic start__shifter_right_tc__width_1024__shift_0__pad_0;

logic start__shifter_right_tc__width_1024__shift_1__pad_0;

logic start__shifter_right_tc__width_1024__shift_2__pad_0;

logic start__shifter_right_tc__width_1024__shift_3__pad_0;

logic start__shifter_right_tc__width_1024__shift_4__pad_0;

logic start__shifter_right_tc__width_1024__shift_5__pad_0;

logic start__shifter_right_tc__width_1024__shift_6__pad_0;

logic start__shifter_right_tc__width_1024__shift_7__pad_0;

logic start__shifter_right_tc__width_1024__shift_512__pad_0;

logic start__shifter_right_tc__width_1024__shift_1023__pad_0;

logic start__shifter_right_tc__width_1024__shift_1024__pad_0;

logic start__shifter_right_tc__width_1024__shift_1025__pad_0;

logic start__shifter_right_tc__width_1024__shift_1536__pad_0;

logic start__shifter_right_tc__width_1024__shift_2047__pad_0;

logic start__shifter_right_tc__width_1024__shift_2048__pad_0;

logic start__shifter_right_tc__width_1024__shift_0__pad_1;

logic start__shifter_right_tc__width_1024__shift_1__pad_1;

logic start__shifter_right_tc__width_1024__shift_2__pad_1;

logic start__shifter_right_tc__width_1024__shift_3__pad_1;

logic start__shifter_right_tc__width_1024__shift_4__pad_1;

logic start__shifter_right_tc__width_1024__shift_5__pad_1;

logic start__shifter_right_tc__width_1024__shift_6__pad_1;

logic start__shifter_right_tc__width_1024__shift_7__pad_1;

logic start__shifter_right_tc__width_1024__shift_512__pad_1;

logic start__shifter_right_tc__width_1024__shift_1023__pad_1;

logic start__shifter_right_tc__width_1024__shift_1024__pad_1;

logic start__shifter_right_tc__width_1024__shift_1025__pad_1;

logic start__shifter_right_tc__width_1024__shift_1536__pad_1;

logic start__shifter_right_tc__width_1024__shift_2047__pad_1;

logic start__shifter_right_tc__width_1024__shift_2048__pad_1;



shifter_right_tc #(.WIDTH(1), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_1__shift_0__pad_0 (.start(start__shifter_right_tc__width_1__shift_0__pad_0));

shifter_right_tc #(.WIDTH(1), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_1__shift_1__pad_0 (.start(start__shifter_right_tc__width_1__shift_1__pad_0));

shifter_right_tc #(.WIDTH(1), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_1__shift_0__pad_1 (.start(start__shifter_right_tc__width_1__shift_0__pad_1));

shifter_right_tc #(.WIDTH(1), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_1__shift_1__pad_1 (.start(start__shifter_right_tc__width_1__shift_1__pad_1));

shifter_right_tc #(.WIDTH(2), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_2__shift_0__pad_0 (.start(start__shifter_right_tc__width_2__shift_0__pad_0));

shifter_right_tc #(.WIDTH(2), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_2__shift_1__pad_0 (.start(start__shifter_right_tc__width_2__shift_1__pad_0));

shifter_right_tc #(.WIDTH(2), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_2__shift_2__pad_0 (.start(start__shifter_right_tc__width_2__shift_2__pad_0));

shifter_right_tc #(.WIDTH(2), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_2__shift_3__pad_0 (.start(start__shifter_right_tc__width_2__shift_3__pad_0));

shifter_right_tc #(.WIDTH(2), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_2__shift_0__pad_1 (.start(start__shifter_right_tc__width_2__shift_0__pad_1));

shifter_right_tc #(.WIDTH(2), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_2__shift_1__pad_1 (.start(start__shifter_right_tc__width_2__shift_1__pad_1));

shifter_right_tc #(.WIDTH(2), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_2__shift_2__pad_1 (.start(start__shifter_right_tc__width_2__shift_2__pad_1));

shifter_right_tc #(.WIDTH(2), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_2__shift_3__pad_1 (.start(start__shifter_right_tc__width_2__shift_3__pad_1));

shifter_right_tc #(.WIDTH(3), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_3__shift_0__pad_0 (.start(start__shifter_right_tc__width_3__shift_0__pad_0));

shifter_right_tc #(.WIDTH(3), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_3__shift_1__pad_0 (.start(start__shifter_right_tc__width_3__shift_1__pad_0));

shifter_right_tc #(.WIDTH(3), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_3__shift_2__pad_0 (.start(start__shifter_right_tc__width_3__shift_2__pad_0));

shifter_right_tc #(.WIDTH(3), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_3__shift_3__pad_0 (.start(start__shifter_right_tc__width_3__shift_3__pad_0));

shifter_right_tc #(.WIDTH(3), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_3__shift_4__pad_0 (.start(start__shifter_right_tc__width_3__shift_4__pad_0));

shifter_right_tc #(.WIDTH(3), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_3__shift_5__pad_0 (.start(start__shifter_right_tc__width_3__shift_5__pad_0));

shifter_right_tc #(.WIDTH(3), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_3__shift_0__pad_1 (.start(start__shifter_right_tc__width_3__shift_0__pad_1));

shifter_right_tc #(.WIDTH(3), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_3__shift_1__pad_1 (.start(start__shifter_right_tc__width_3__shift_1__pad_1));

shifter_right_tc #(.WIDTH(3), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_3__shift_2__pad_1 (.start(start__shifter_right_tc__width_3__shift_2__pad_1));

shifter_right_tc #(.WIDTH(3), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_3__shift_3__pad_1 (.start(start__shifter_right_tc__width_3__shift_3__pad_1));

shifter_right_tc #(.WIDTH(3), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_3__shift_4__pad_1 (.start(start__shifter_right_tc__width_3__shift_4__pad_1));

shifter_right_tc #(.WIDTH(3), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_3__shift_5__pad_1 (.start(start__shifter_right_tc__width_3__shift_5__pad_1));

shifter_right_tc #(.WIDTH(4), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_4__shift_0__pad_0 (.start(start__shifter_right_tc__width_4__shift_0__pad_0));

shifter_right_tc #(.WIDTH(4), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_4__shift_1__pad_0 (.start(start__shifter_right_tc__width_4__shift_1__pad_0));

shifter_right_tc #(.WIDTH(4), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_4__shift_2__pad_0 (.start(start__shifter_right_tc__width_4__shift_2__pad_0));

shifter_right_tc #(.WIDTH(4), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_4__shift_3__pad_0 (.start(start__shifter_right_tc__width_4__shift_3__pad_0));

shifter_right_tc #(.WIDTH(4), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_4__shift_4__pad_0 (.start(start__shifter_right_tc__width_4__shift_4__pad_0));

shifter_right_tc #(.WIDTH(4), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_4__shift_5__pad_0 (.start(start__shifter_right_tc__width_4__shift_5__pad_0));

shifter_right_tc #(.WIDTH(4), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_4__shift_6__pad_0 (.start(start__shifter_right_tc__width_4__shift_6__pad_0));

shifter_right_tc #(.WIDTH(4), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_4__shift_7__pad_0 (.start(start__shifter_right_tc__width_4__shift_7__pad_0));

shifter_right_tc #(.WIDTH(4), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_4__shift_0__pad_1 (.start(start__shifter_right_tc__width_4__shift_0__pad_1));

shifter_right_tc #(.WIDTH(4), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_4__shift_1__pad_1 (.start(start__shifter_right_tc__width_4__shift_1__pad_1));

shifter_right_tc #(.WIDTH(4), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_4__shift_2__pad_1 (.start(start__shifter_right_tc__width_4__shift_2__pad_1));

shifter_right_tc #(.WIDTH(4), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_4__shift_3__pad_1 (.start(start__shifter_right_tc__width_4__shift_3__pad_1));

shifter_right_tc #(.WIDTH(4), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_4__shift_4__pad_1 (.start(start__shifter_right_tc__width_4__shift_4__pad_1));

shifter_right_tc #(.WIDTH(4), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_4__shift_5__pad_1 (.start(start__shifter_right_tc__width_4__shift_5__pad_1));

shifter_right_tc #(.WIDTH(4), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_4__shift_6__pad_1 (.start(start__shifter_right_tc__width_4__shift_6__pad_1));

shifter_right_tc #(.WIDTH(4), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_4__shift_7__pad_1 (.start(start__shifter_right_tc__width_4__shift_7__pad_1));

shifter_right_tc #(.WIDTH(5), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_5__shift_0__pad_0 (.start(start__shifter_right_tc__width_5__shift_0__pad_0));

shifter_right_tc #(.WIDTH(5), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_5__shift_1__pad_0 (.start(start__shifter_right_tc__width_5__shift_1__pad_0));

shifter_right_tc #(.WIDTH(5), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_5__shift_2__pad_0 (.start(start__shifter_right_tc__width_5__shift_2__pad_0));

shifter_right_tc #(.WIDTH(5), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_5__shift_3__pad_0 (.start(start__shifter_right_tc__width_5__shift_3__pad_0));

shifter_right_tc #(.WIDTH(5), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_5__shift_4__pad_0 (.start(start__shifter_right_tc__width_5__shift_4__pad_0));

shifter_right_tc #(.WIDTH(5), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_5__shift_5__pad_0 (.start(start__shifter_right_tc__width_5__shift_5__pad_0));

shifter_right_tc #(.WIDTH(5), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_5__shift_6__pad_0 (.start(start__shifter_right_tc__width_5__shift_6__pad_0));

shifter_right_tc #(.WIDTH(5), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_5__shift_7__pad_0 (.start(start__shifter_right_tc__width_5__shift_7__pad_0));

shifter_right_tc #(.WIDTH(5), .SHIFT(8), .PAD_VALUE(0)) shifter_right_tc__width_5__shift_8__pad_0 (.start(start__shifter_right_tc__width_5__shift_8__pad_0));

shifter_right_tc #(.WIDTH(5), .SHIFT(9), .PAD_VALUE(0)) shifter_right_tc__width_5__shift_9__pad_0 (.start(start__shifter_right_tc__width_5__shift_9__pad_0));

shifter_right_tc #(.WIDTH(5), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_5__shift_0__pad_1 (.start(start__shifter_right_tc__width_5__shift_0__pad_1));

shifter_right_tc #(.WIDTH(5), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_5__shift_1__pad_1 (.start(start__shifter_right_tc__width_5__shift_1__pad_1));

shifter_right_tc #(.WIDTH(5), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_5__shift_2__pad_1 (.start(start__shifter_right_tc__width_5__shift_2__pad_1));

shifter_right_tc #(.WIDTH(5), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_5__shift_3__pad_1 (.start(start__shifter_right_tc__width_5__shift_3__pad_1));

shifter_right_tc #(.WIDTH(5), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_5__shift_4__pad_1 (.start(start__shifter_right_tc__width_5__shift_4__pad_1));

shifter_right_tc #(.WIDTH(5), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_5__shift_5__pad_1 (.start(start__shifter_right_tc__width_5__shift_5__pad_1));

shifter_right_tc #(.WIDTH(5), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_5__shift_6__pad_1 (.start(start__shifter_right_tc__width_5__shift_6__pad_1));

shifter_right_tc #(.WIDTH(5), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_5__shift_7__pad_1 (.start(start__shifter_right_tc__width_5__shift_7__pad_1));

shifter_right_tc #(.WIDTH(5), .SHIFT(8), .PAD_VALUE(1)) shifter_right_tc__width_5__shift_8__pad_1 (.start(start__shifter_right_tc__width_5__shift_8__pad_1));

shifter_right_tc #(.WIDTH(5), .SHIFT(9), .PAD_VALUE(1)) shifter_right_tc__width_5__shift_9__pad_1 (.start(start__shifter_right_tc__width_5__shift_9__pad_1));

shifter_right_tc #(.WIDTH(6), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_6__shift_0__pad_0 (.start(start__shifter_right_tc__width_6__shift_0__pad_0));

shifter_right_tc #(.WIDTH(6), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_6__shift_1__pad_0 (.start(start__shifter_right_tc__width_6__shift_1__pad_0));

shifter_right_tc #(.WIDTH(6), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_6__shift_2__pad_0 (.start(start__shifter_right_tc__width_6__shift_2__pad_0));

shifter_right_tc #(.WIDTH(6), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_6__shift_3__pad_0 (.start(start__shifter_right_tc__width_6__shift_3__pad_0));

shifter_right_tc #(.WIDTH(6), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_6__shift_4__pad_0 (.start(start__shifter_right_tc__width_6__shift_4__pad_0));

shifter_right_tc #(.WIDTH(6), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_6__shift_5__pad_0 (.start(start__shifter_right_tc__width_6__shift_5__pad_0));

shifter_right_tc #(.WIDTH(6), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_6__shift_6__pad_0 (.start(start__shifter_right_tc__width_6__shift_6__pad_0));

shifter_right_tc #(.WIDTH(6), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_6__shift_7__pad_0 (.start(start__shifter_right_tc__width_6__shift_7__pad_0));

shifter_right_tc #(.WIDTH(6), .SHIFT(8), .PAD_VALUE(0)) shifter_right_tc__width_6__shift_8__pad_0 (.start(start__shifter_right_tc__width_6__shift_8__pad_0));

shifter_right_tc #(.WIDTH(6), .SHIFT(9), .PAD_VALUE(0)) shifter_right_tc__width_6__shift_9__pad_0 (.start(start__shifter_right_tc__width_6__shift_9__pad_0));

shifter_right_tc #(.WIDTH(6), .SHIFT(10), .PAD_VALUE(0)) shifter_right_tc__width_6__shift_10__pad_0 (.start(start__shifter_right_tc__width_6__shift_10__pad_0));

shifter_right_tc #(.WIDTH(6), .SHIFT(11), .PAD_VALUE(0)) shifter_right_tc__width_6__shift_11__pad_0 (.start(start__shifter_right_tc__width_6__shift_11__pad_0));

shifter_right_tc #(.WIDTH(6), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_6__shift_0__pad_1 (.start(start__shifter_right_tc__width_6__shift_0__pad_1));

shifter_right_tc #(.WIDTH(6), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_6__shift_1__pad_1 (.start(start__shifter_right_tc__width_6__shift_1__pad_1));

shifter_right_tc #(.WIDTH(6), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_6__shift_2__pad_1 (.start(start__shifter_right_tc__width_6__shift_2__pad_1));

shifter_right_tc #(.WIDTH(6), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_6__shift_3__pad_1 (.start(start__shifter_right_tc__width_6__shift_3__pad_1));

shifter_right_tc #(.WIDTH(6), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_6__shift_4__pad_1 (.start(start__shifter_right_tc__width_6__shift_4__pad_1));

shifter_right_tc #(.WIDTH(6), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_6__shift_5__pad_1 (.start(start__shifter_right_tc__width_6__shift_5__pad_1));

shifter_right_tc #(.WIDTH(6), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_6__shift_6__pad_1 (.start(start__shifter_right_tc__width_6__shift_6__pad_1));

shifter_right_tc #(.WIDTH(6), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_6__shift_7__pad_1 (.start(start__shifter_right_tc__width_6__shift_7__pad_1));

shifter_right_tc #(.WIDTH(6), .SHIFT(8), .PAD_VALUE(1)) shifter_right_tc__width_6__shift_8__pad_1 (.start(start__shifter_right_tc__width_6__shift_8__pad_1));

shifter_right_tc #(.WIDTH(6), .SHIFT(9), .PAD_VALUE(1)) shifter_right_tc__width_6__shift_9__pad_1 (.start(start__shifter_right_tc__width_6__shift_9__pad_1));

shifter_right_tc #(.WIDTH(6), .SHIFT(10), .PAD_VALUE(1)) shifter_right_tc__width_6__shift_10__pad_1 (.start(start__shifter_right_tc__width_6__shift_10__pad_1));

shifter_right_tc #(.WIDTH(6), .SHIFT(11), .PAD_VALUE(1)) shifter_right_tc__width_6__shift_11__pad_1 (.start(start__shifter_right_tc__width_6__shift_11__pad_1));

shifter_right_tc #(.WIDTH(7), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_7__shift_0__pad_0 (.start(start__shifter_right_tc__width_7__shift_0__pad_0));

shifter_right_tc #(.WIDTH(7), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_7__shift_1__pad_0 (.start(start__shifter_right_tc__width_7__shift_1__pad_0));

shifter_right_tc #(.WIDTH(7), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_7__shift_2__pad_0 (.start(start__shifter_right_tc__width_7__shift_2__pad_0));

shifter_right_tc #(.WIDTH(7), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_7__shift_3__pad_0 (.start(start__shifter_right_tc__width_7__shift_3__pad_0));

shifter_right_tc #(.WIDTH(7), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_7__shift_4__pad_0 (.start(start__shifter_right_tc__width_7__shift_4__pad_0));

shifter_right_tc #(.WIDTH(7), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_7__shift_5__pad_0 (.start(start__shifter_right_tc__width_7__shift_5__pad_0));

shifter_right_tc #(.WIDTH(7), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_7__shift_6__pad_0 (.start(start__shifter_right_tc__width_7__shift_6__pad_0));

shifter_right_tc #(.WIDTH(7), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_7__shift_7__pad_0 (.start(start__shifter_right_tc__width_7__shift_7__pad_0));

shifter_right_tc #(.WIDTH(7), .SHIFT(8), .PAD_VALUE(0)) shifter_right_tc__width_7__shift_8__pad_0 (.start(start__shifter_right_tc__width_7__shift_8__pad_0));

shifter_right_tc #(.WIDTH(7), .SHIFT(9), .PAD_VALUE(0)) shifter_right_tc__width_7__shift_9__pad_0 (.start(start__shifter_right_tc__width_7__shift_9__pad_0));

shifter_right_tc #(.WIDTH(7), .SHIFT(10), .PAD_VALUE(0)) shifter_right_tc__width_7__shift_10__pad_0 (.start(start__shifter_right_tc__width_7__shift_10__pad_0));

shifter_right_tc #(.WIDTH(7), .SHIFT(11), .PAD_VALUE(0)) shifter_right_tc__width_7__shift_11__pad_0 (.start(start__shifter_right_tc__width_7__shift_11__pad_0));

shifter_right_tc #(.WIDTH(7), .SHIFT(12), .PAD_VALUE(0)) shifter_right_tc__width_7__shift_12__pad_0 (.start(start__shifter_right_tc__width_7__shift_12__pad_0));

shifter_right_tc #(.WIDTH(7), .SHIFT(13), .PAD_VALUE(0)) shifter_right_tc__width_7__shift_13__pad_0 (.start(start__shifter_right_tc__width_7__shift_13__pad_0));

shifter_right_tc #(.WIDTH(7), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_7__shift_0__pad_1 (.start(start__shifter_right_tc__width_7__shift_0__pad_1));

shifter_right_tc #(.WIDTH(7), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_7__shift_1__pad_1 (.start(start__shifter_right_tc__width_7__shift_1__pad_1));

shifter_right_tc #(.WIDTH(7), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_7__shift_2__pad_1 (.start(start__shifter_right_tc__width_7__shift_2__pad_1));

shifter_right_tc #(.WIDTH(7), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_7__shift_3__pad_1 (.start(start__shifter_right_tc__width_7__shift_3__pad_1));

shifter_right_tc #(.WIDTH(7), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_7__shift_4__pad_1 (.start(start__shifter_right_tc__width_7__shift_4__pad_1));

shifter_right_tc #(.WIDTH(7), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_7__shift_5__pad_1 (.start(start__shifter_right_tc__width_7__shift_5__pad_1));

shifter_right_tc #(.WIDTH(7), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_7__shift_6__pad_1 (.start(start__shifter_right_tc__width_7__shift_6__pad_1));

shifter_right_tc #(.WIDTH(7), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_7__shift_7__pad_1 (.start(start__shifter_right_tc__width_7__shift_7__pad_1));

shifter_right_tc #(.WIDTH(7), .SHIFT(8), .PAD_VALUE(1)) shifter_right_tc__width_7__shift_8__pad_1 (.start(start__shifter_right_tc__width_7__shift_8__pad_1));

shifter_right_tc #(.WIDTH(7), .SHIFT(9), .PAD_VALUE(1)) shifter_right_tc__width_7__shift_9__pad_1 (.start(start__shifter_right_tc__width_7__shift_9__pad_1));

shifter_right_tc #(.WIDTH(7), .SHIFT(10), .PAD_VALUE(1)) shifter_right_tc__width_7__shift_10__pad_1 (.start(start__shifter_right_tc__width_7__shift_10__pad_1));

shifter_right_tc #(.WIDTH(7), .SHIFT(11), .PAD_VALUE(1)) shifter_right_tc__width_7__shift_11__pad_1 (.start(start__shifter_right_tc__width_7__shift_11__pad_1));

shifter_right_tc #(.WIDTH(7), .SHIFT(12), .PAD_VALUE(1)) shifter_right_tc__width_7__shift_12__pad_1 (.start(start__shifter_right_tc__width_7__shift_12__pad_1));

shifter_right_tc #(.WIDTH(7), .SHIFT(13), .PAD_VALUE(1)) shifter_right_tc__width_7__shift_13__pad_1 (.start(start__shifter_right_tc__width_7__shift_13__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_0__pad_0 (.start(start__shifter_right_tc__width_8__shift_0__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_1__pad_0 (.start(start__shifter_right_tc__width_8__shift_1__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_2__pad_0 (.start(start__shifter_right_tc__width_8__shift_2__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_3__pad_0 (.start(start__shifter_right_tc__width_8__shift_3__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_4__pad_0 (.start(start__shifter_right_tc__width_8__shift_4__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_5__pad_0 (.start(start__shifter_right_tc__width_8__shift_5__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_6__pad_0 (.start(start__shifter_right_tc__width_8__shift_6__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_7__pad_0 (.start(start__shifter_right_tc__width_8__shift_7__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(8), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_8__pad_0 (.start(start__shifter_right_tc__width_8__shift_8__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(9), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_9__pad_0 (.start(start__shifter_right_tc__width_8__shift_9__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(10), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_10__pad_0 (.start(start__shifter_right_tc__width_8__shift_10__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(11), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_11__pad_0 (.start(start__shifter_right_tc__width_8__shift_11__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(12), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_12__pad_0 (.start(start__shifter_right_tc__width_8__shift_12__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(13), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_13__pad_0 (.start(start__shifter_right_tc__width_8__shift_13__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(14), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_14__pad_0 (.start(start__shifter_right_tc__width_8__shift_14__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(15), .PAD_VALUE(0)) shifter_right_tc__width_8__shift_15__pad_0 (.start(start__shifter_right_tc__width_8__shift_15__pad_0));

shifter_right_tc #(.WIDTH(8), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_0__pad_1 (.start(start__shifter_right_tc__width_8__shift_0__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_1__pad_1 (.start(start__shifter_right_tc__width_8__shift_1__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_2__pad_1 (.start(start__shifter_right_tc__width_8__shift_2__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_3__pad_1 (.start(start__shifter_right_tc__width_8__shift_3__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_4__pad_1 (.start(start__shifter_right_tc__width_8__shift_4__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_5__pad_1 (.start(start__shifter_right_tc__width_8__shift_5__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_6__pad_1 (.start(start__shifter_right_tc__width_8__shift_6__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_7__pad_1 (.start(start__shifter_right_tc__width_8__shift_7__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(8), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_8__pad_1 (.start(start__shifter_right_tc__width_8__shift_8__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(9), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_9__pad_1 (.start(start__shifter_right_tc__width_8__shift_9__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(10), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_10__pad_1 (.start(start__shifter_right_tc__width_8__shift_10__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(11), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_11__pad_1 (.start(start__shifter_right_tc__width_8__shift_11__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(12), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_12__pad_1 (.start(start__shifter_right_tc__width_8__shift_12__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(13), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_13__pad_1 (.start(start__shifter_right_tc__width_8__shift_13__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(14), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_14__pad_1 (.start(start__shifter_right_tc__width_8__shift_14__pad_1));

shifter_right_tc #(.WIDTH(8), .SHIFT(15), .PAD_VALUE(1)) shifter_right_tc__width_8__shift_15__pad_1 (.start(start__shifter_right_tc__width_8__shift_15__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_0__pad_0 (.start(start__shifter_right_tc__width_9__shift_0__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_1__pad_0 (.start(start__shifter_right_tc__width_9__shift_1__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_2__pad_0 (.start(start__shifter_right_tc__width_9__shift_2__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_3__pad_0 (.start(start__shifter_right_tc__width_9__shift_3__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_4__pad_0 (.start(start__shifter_right_tc__width_9__shift_4__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_5__pad_0 (.start(start__shifter_right_tc__width_9__shift_5__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_6__pad_0 (.start(start__shifter_right_tc__width_9__shift_6__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_7__pad_0 (.start(start__shifter_right_tc__width_9__shift_7__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(8), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_8__pad_0 (.start(start__shifter_right_tc__width_9__shift_8__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(9), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_9__pad_0 (.start(start__shifter_right_tc__width_9__shift_9__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(10), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_10__pad_0 (.start(start__shifter_right_tc__width_9__shift_10__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(11), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_11__pad_0 (.start(start__shifter_right_tc__width_9__shift_11__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(12), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_12__pad_0 (.start(start__shifter_right_tc__width_9__shift_12__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(13), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_13__pad_0 (.start(start__shifter_right_tc__width_9__shift_13__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(14), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_14__pad_0 (.start(start__shifter_right_tc__width_9__shift_14__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(15), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_15__pad_0 (.start(start__shifter_right_tc__width_9__shift_15__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(16), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_16__pad_0 (.start(start__shifter_right_tc__width_9__shift_16__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(17), .PAD_VALUE(0)) shifter_right_tc__width_9__shift_17__pad_0 (.start(start__shifter_right_tc__width_9__shift_17__pad_0));

shifter_right_tc #(.WIDTH(9), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_0__pad_1 (.start(start__shifter_right_tc__width_9__shift_0__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_1__pad_1 (.start(start__shifter_right_tc__width_9__shift_1__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_2__pad_1 (.start(start__shifter_right_tc__width_9__shift_2__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_3__pad_1 (.start(start__shifter_right_tc__width_9__shift_3__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_4__pad_1 (.start(start__shifter_right_tc__width_9__shift_4__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_5__pad_1 (.start(start__shifter_right_tc__width_9__shift_5__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_6__pad_1 (.start(start__shifter_right_tc__width_9__shift_6__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_7__pad_1 (.start(start__shifter_right_tc__width_9__shift_7__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(8), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_8__pad_1 (.start(start__shifter_right_tc__width_9__shift_8__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(9), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_9__pad_1 (.start(start__shifter_right_tc__width_9__shift_9__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(10), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_10__pad_1 (.start(start__shifter_right_tc__width_9__shift_10__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(11), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_11__pad_1 (.start(start__shifter_right_tc__width_9__shift_11__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(12), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_12__pad_1 (.start(start__shifter_right_tc__width_9__shift_12__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(13), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_13__pad_1 (.start(start__shifter_right_tc__width_9__shift_13__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(14), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_14__pad_1 (.start(start__shifter_right_tc__width_9__shift_14__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(15), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_15__pad_1 (.start(start__shifter_right_tc__width_9__shift_15__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(16), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_16__pad_1 (.start(start__shifter_right_tc__width_9__shift_16__pad_1));

shifter_right_tc #(.WIDTH(9), .SHIFT(17), .PAD_VALUE(1)) shifter_right_tc__width_9__shift_17__pad_1 (.start(start__shifter_right_tc__width_9__shift_17__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_0__pad_0 (.start(start__shifter_right_tc__width_10__shift_0__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_1__pad_0 (.start(start__shifter_right_tc__width_10__shift_1__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_2__pad_0 (.start(start__shifter_right_tc__width_10__shift_2__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_3__pad_0 (.start(start__shifter_right_tc__width_10__shift_3__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_4__pad_0 (.start(start__shifter_right_tc__width_10__shift_4__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_5__pad_0 (.start(start__shifter_right_tc__width_10__shift_5__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_6__pad_0 (.start(start__shifter_right_tc__width_10__shift_6__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_7__pad_0 (.start(start__shifter_right_tc__width_10__shift_7__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(8), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_8__pad_0 (.start(start__shifter_right_tc__width_10__shift_8__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(9), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_9__pad_0 (.start(start__shifter_right_tc__width_10__shift_9__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(10), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_10__pad_0 (.start(start__shifter_right_tc__width_10__shift_10__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(11), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_11__pad_0 (.start(start__shifter_right_tc__width_10__shift_11__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(12), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_12__pad_0 (.start(start__shifter_right_tc__width_10__shift_12__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(13), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_13__pad_0 (.start(start__shifter_right_tc__width_10__shift_13__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(14), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_14__pad_0 (.start(start__shifter_right_tc__width_10__shift_14__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(15), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_15__pad_0 (.start(start__shifter_right_tc__width_10__shift_15__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(16), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_16__pad_0 (.start(start__shifter_right_tc__width_10__shift_16__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(17), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_17__pad_0 (.start(start__shifter_right_tc__width_10__shift_17__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(18), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_18__pad_0 (.start(start__shifter_right_tc__width_10__shift_18__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(19), .PAD_VALUE(0)) shifter_right_tc__width_10__shift_19__pad_0 (.start(start__shifter_right_tc__width_10__shift_19__pad_0));

shifter_right_tc #(.WIDTH(10), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_0__pad_1 (.start(start__shifter_right_tc__width_10__shift_0__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_1__pad_1 (.start(start__shifter_right_tc__width_10__shift_1__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_2__pad_1 (.start(start__shifter_right_tc__width_10__shift_2__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_3__pad_1 (.start(start__shifter_right_tc__width_10__shift_3__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_4__pad_1 (.start(start__shifter_right_tc__width_10__shift_4__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_5__pad_1 (.start(start__shifter_right_tc__width_10__shift_5__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_6__pad_1 (.start(start__shifter_right_tc__width_10__shift_6__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_7__pad_1 (.start(start__shifter_right_tc__width_10__shift_7__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(8), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_8__pad_1 (.start(start__shifter_right_tc__width_10__shift_8__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(9), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_9__pad_1 (.start(start__shifter_right_tc__width_10__shift_9__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(10), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_10__pad_1 (.start(start__shifter_right_tc__width_10__shift_10__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(11), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_11__pad_1 (.start(start__shifter_right_tc__width_10__shift_11__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(12), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_12__pad_1 (.start(start__shifter_right_tc__width_10__shift_12__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(13), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_13__pad_1 (.start(start__shifter_right_tc__width_10__shift_13__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(14), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_14__pad_1 (.start(start__shifter_right_tc__width_10__shift_14__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(15), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_15__pad_1 (.start(start__shifter_right_tc__width_10__shift_15__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(16), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_16__pad_1 (.start(start__shifter_right_tc__width_10__shift_16__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(17), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_17__pad_1 (.start(start__shifter_right_tc__width_10__shift_17__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(18), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_18__pad_1 (.start(start__shifter_right_tc__width_10__shift_18__pad_1));

shifter_right_tc #(.WIDTH(10), .SHIFT(19), .PAD_VALUE(1)) shifter_right_tc__width_10__shift_19__pad_1 (.start(start__shifter_right_tc__width_10__shift_19__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_0__pad_0 (.start(start__shifter_right_tc__width_11__shift_0__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_1__pad_0 (.start(start__shifter_right_tc__width_11__shift_1__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_2__pad_0 (.start(start__shifter_right_tc__width_11__shift_2__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_3__pad_0 (.start(start__shifter_right_tc__width_11__shift_3__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_4__pad_0 (.start(start__shifter_right_tc__width_11__shift_4__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_5__pad_0 (.start(start__shifter_right_tc__width_11__shift_5__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_6__pad_0 (.start(start__shifter_right_tc__width_11__shift_6__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_7__pad_0 (.start(start__shifter_right_tc__width_11__shift_7__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(8), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_8__pad_0 (.start(start__shifter_right_tc__width_11__shift_8__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(9), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_9__pad_0 (.start(start__shifter_right_tc__width_11__shift_9__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(10), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_10__pad_0 (.start(start__shifter_right_tc__width_11__shift_10__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(11), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_11__pad_0 (.start(start__shifter_right_tc__width_11__shift_11__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(12), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_12__pad_0 (.start(start__shifter_right_tc__width_11__shift_12__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(13), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_13__pad_0 (.start(start__shifter_right_tc__width_11__shift_13__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(14), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_14__pad_0 (.start(start__shifter_right_tc__width_11__shift_14__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(15), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_15__pad_0 (.start(start__shifter_right_tc__width_11__shift_15__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(16), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_16__pad_0 (.start(start__shifter_right_tc__width_11__shift_16__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(17), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_17__pad_0 (.start(start__shifter_right_tc__width_11__shift_17__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(18), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_18__pad_0 (.start(start__shifter_right_tc__width_11__shift_18__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(19), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_19__pad_0 (.start(start__shifter_right_tc__width_11__shift_19__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(20), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_20__pad_0 (.start(start__shifter_right_tc__width_11__shift_20__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(21), .PAD_VALUE(0)) shifter_right_tc__width_11__shift_21__pad_0 (.start(start__shifter_right_tc__width_11__shift_21__pad_0));

shifter_right_tc #(.WIDTH(11), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_0__pad_1 (.start(start__shifter_right_tc__width_11__shift_0__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_1__pad_1 (.start(start__shifter_right_tc__width_11__shift_1__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_2__pad_1 (.start(start__shifter_right_tc__width_11__shift_2__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_3__pad_1 (.start(start__shifter_right_tc__width_11__shift_3__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_4__pad_1 (.start(start__shifter_right_tc__width_11__shift_4__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_5__pad_1 (.start(start__shifter_right_tc__width_11__shift_5__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_6__pad_1 (.start(start__shifter_right_tc__width_11__shift_6__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_7__pad_1 (.start(start__shifter_right_tc__width_11__shift_7__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(8), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_8__pad_1 (.start(start__shifter_right_tc__width_11__shift_8__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(9), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_9__pad_1 (.start(start__shifter_right_tc__width_11__shift_9__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(10), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_10__pad_1 (.start(start__shifter_right_tc__width_11__shift_10__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(11), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_11__pad_1 (.start(start__shifter_right_tc__width_11__shift_11__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(12), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_12__pad_1 (.start(start__shifter_right_tc__width_11__shift_12__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(13), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_13__pad_1 (.start(start__shifter_right_tc__width_11__shift_13__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(14), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_14__pad_1 (.start(start__shifter_right_tc__width_11__shift_14__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(15), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_15__pad_1 (.start(start__shifter_right_tc__width_11__shift_15__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(16), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_16__pad_1 (.start(start__shifter_right_tc__width_11__shift_16__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(17), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_17__pad_1 (.start(start__shifter_right_tc__width_11__shift_17__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(18), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_18__pad_1 (.start(start__shifter_right_tc__width_11__shift_18__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(19), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_19__pad_1 (.start(start__shifter_right_tc__width_11__shift_19__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(20), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_20__pad_1 (.start(start__shifter_right_tc__width_11__shift_20__pad_1));

shifter_right_tc #(.WIDTH(11), .SHIFT(21), .PAD_VALUE(1)) shifter_right_tc__width_11__shift_21__pad_1 (.start(start__shifter_right_tc__width_11__shift_21__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_0__pad_0 (.start(start__shifter_right_tc__width_12__shift_0__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_1__pad_0 (.start(start__shifter_right_tc__width_12__shift_1__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_2__pad_0 (.start(start__shifter_right_tc__width_12__shift_2__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_3__pad_0 (.start(start__shifter_right_tc__width_12__shift_3__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_4__pad_0 (.start(start__shifter_right_tc__width_12__shift_4__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_5__pad_0 (.start(start__shifter_right_tc__width_12__shift_5__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_6__pad_0 (.start(start__shifter_right_tc__width_12__shift_6__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_7__pad_0 (.start(start__shifter_right_tc__width_12__shift_7__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(8), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_8__pad_0 (.start(start__shifter_right_tc__width_12__shift_8__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(9), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_9__pad_0 (.start(start__shifter_right_tc__width_12__shift_9__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(10), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_10__pad_0 (.start(start__shifter_right_tc__width_12__shift_10__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(11), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_11__pad_0 (.start(start__shifter_right_tc__width_12__shift_11__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(12), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_12__pad_0 (.start(start__shifter_right_tc__width_12__shift_12__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(13), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_13__pad_0 (.start(start__shifter_right_tc__width_12__shift_13__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(14), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_14__pad_0 (.start(start__shifter_right_tc__width_12__shift_14__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(15), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_15__pad_0 (.start(start__shifter_right_tc__width_12__shift_15__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(16), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_16__pad_0 (.start(start__shifter_right_tc__width_12__shift_16__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(17), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_17__pad_0 (.start(start__shifter_right_tc__width_12__shift_17__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(18), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_18__pad_0 (.start(start__shifter_right_tc__width_12__shift_18__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(19), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_19__pad_0 (.start(start__shifter_right_tc__width_12__shift_19__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(20), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_20__pad_0 (.start(start__shifter_right_tc__width_12__shift_20__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(21), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_21__pad_0 (.start(start__shifter_right_tc__width_12__shift_21__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(22), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_22__pad_0 (.start(start__shifter_right_tc__width_12__shift_22__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(23), .PAD_VALUE(0)) shifter_right_tc__width_12__shift_23__pad_0 (.start(start__shifter_right_tc__width_12__shift_23__pad_0));

shifter_right_tc #(.WIDTH(12), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_0__pad_1 (.start(start__shifter_right_tc__width_12__shift_0__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_1__pad_1 (.start(start__shifter_right_tc__width_12__shift_1__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_2__pad_1 (.start(start__shifter_right_tc__width_12__shift_2__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_3__pad_1 (.start(start__shifter_right_tc__width_12__shift_3__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_4__pad_1 (.start(start__shifter_right_tc__width_12__shift_4__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_5__pad_1 (.start(start__shifter_right_tc__width_12__shift_5__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_6__pad_1 (.start(start__shifter_right_tc__width_12__shift_6__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_7__pad_1 (.start(start__shifter_right_tc__width_12__shift_7__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(8), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_8__pad_1 (.start(start__shifter_right_tc__width_12__shift_8__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(9), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_9__pad_1 (.start(start__shifter_right_tc__width_12__shift_9__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(10), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_10__pad_1 (.start(start__shifter_right_tc__width_12__shift_10__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(11), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_11__pad_1 (.start(start__shifter_right_tc__width_12__shift_11__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(12), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_12__pad_1 (.start(start__shifter_right_tc__width_12__shift_12__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(13), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_13__pad_1 (.start(start__shifter_right_tc__width_12__shift_13__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(14), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_14__pad_1 (.start(start__shifter_right_tc__width_12__shift_14__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(15), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_15__pad_1 (.start(start__shifter_right_tc__width_12__shift_15__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(16), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_16__pad_1 (.start(start__shifter_right_tc__width_12__shift_16__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(17), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_17__pad_1 (.start(start__shifter_right_tc__width_12__shift_17__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(18), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_18__pad_1 (.start(start__shifter_right_tc__width_12__shift_18__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(19), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_19__pad_1 (.start(start__shifter_right_tc__width_12__shift_19__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(20), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_20__pad_1 (.start(start__shifter_right_tc__width_12__shift_20__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(21), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_21__pad_1 (.start(start__shifter_right_tc__width_12__shift_21__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(22), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_22__pad_1 (.start(start__shifter_right_tc__width_12__shift_22__pad_1));

shifter_right_tc #(.WIDTH(12), .SHIFT(23), .PAD_VALUE(1)) shifter_right_tc__width_12__shift_23__pad_1 (.start(start__shifter_right_tc__width_12__shift_23__pad_1));

shifter_right_tc #(.WIDTH(16), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_16__shift_0__pad_0 (.start(start__shifter_right_tc__width_16__shift_0__pad_0));

shifter_right_tc #(.WIDTH(16), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_16__shift_1__pad_0 (.start(start__shifter_right_tc__width_16__shift_1__pad_0));

shifter_right_tc #(.WIDTH(16), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_16__shift_2__pad_0 (.start(start__shifter_right_tc__width_16__shift_2__pad_0));

shifter_right_tc #(.WIDTH(16), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_16__shift_3__pad_0 (.start(start__shifter_right_tc__width_16__shift_3__pad_0));

shifter_right_tc #(.WIDTH(16), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_16__shift_4__pad_0 (.start(start__shifter_right_tc__width_16__shift_4__pad_0));

shifter_right_tc #(.WIDTH(16), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_16__shift_5__pad_0 (.start(start__shifter_right_tc__width_16__shift_5__pad_0));

shifter_right_tc #(.WIDTH(16), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_16__shift_6__pad_0 (.start(start__shifter_right_tc__width_16__shift_6__pad_0));

shifter_right_tc #(.WIDTH(16), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_16__shift_7__pad_0 (.start(start__shifter_right_tc__width_16__shift_7__pad_0));

shifter_right_tc #(.WIDTH(16), .SHIFT(8), .PAD_VALUE(0)) shifter_right_tc__width_16__shift_8__pad_0 (.start(start__shifter_right_tc__width_16__shift_8__pad_0));

shifter_right_tc #(.WIDTH(16), .SHIFT(15), .PAD_VALUE(0)) shifter_right_tc__width_16__shift_15__pad_0 (.start(start__shifter_right_tc__width_16__shift_15__pad_0));

shifter_right_tc #(.WIDTH(16), .SHIFT(16), .PAD_VALUE(0)) shifter_right_tc__width_16__shift_16__pad_0 (.start(start__shifter_right_tc__width_16__shift_16__pad_0));

shifter_right_tc #(.WIDTH(16), .SHIFT(17), .PAD_VALUE(0)) shifter_right_tc__width_16__shift_17__pad_0 (.start(start__shifter_right_tc__width_16__shift_17__pad_0));

shifter_right_tc #(.WIDTH(16), .SHIFT(24), .PAD_VALUE(0)) shifter_right_tc__width_16__shift_24__pad_0 (.start(start__shifter_right_tc__width_16__shift_24__pad_0));

shifter_right_tc #(.WIDTH(16), .SHIFT(31), .PAD_VALUE(0)) shifter_right_tc__width_16__shift_31__pad_0 (.start(start__shifter_right_tc__width_16__shift_31__pad_0));

shifter_right_tc #(.WIDTH(16), .SHIFT(32), .PAD_VALUE(0)) shifter_right_tc__width_16__shift_32__pad_0 (.start(start__shifter_right_tc__width_16__shift_32__pad_0));

shifter_right_tc #(.WIDTH(16), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_16__shift_0__pad_1 (.start(start__shifter_right_tc__width_16__shift_0__pad_1));

shifter_right_tc #(.WIDTH(16), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_16__shift_1__pad_1 (.start(start__shifter_right_tc__width_16__shift_1__pad_1));

shifter_right_tc #(.WIDTH(16), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_16__shift_2__pad_1 (.start(start__shifter_right_tc__width_16__shift_2__pad_1));

shifter_right_tc #(.WIDTH(16), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_16__shift_3__pad_1 (.start(start__shifter_right_tc__width_16__shift_3__pad_1));

shifter_right_tc #(.WIDTH(16), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_16__shift_4__pad_1 (.start(start__shifter_right_tc__width_16__shift_4__pad_1));

shifter_right_tc #(.WIDTH(16), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_16__shift_5__pad_1 (.start(start__shifter_right_tc__width_16__shift_5__pad_1));

shifter_right_tc #(.WIDTH(16), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_16__shift_6__pad_1 (.start(start__shifter_right_tc__width_16__shift_6__pad_1));

shifter_right_tc #(.WIDTH(16), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_16__shift_7__pad_1 (.start(start__shifter_right_tc__width_16__shift_7__pad_1));

shifter_right_tc #(.WIDTH(16), .SHIFT(8), .PAD_VALUE(1)) shifter_right_tc__width_16__shift_8__pad_1 (.start(start__shifter_right_tc__width_16__shift_8__pad_1));

shifter_right_tc #(.WIDTH(16), .SHIFT(15), .PAD_VALUE(1)) shifter_right_tc__width_16__shift_15__pad_1 (.start(start__shifter_right_tc__width_16__shift_15__pad_1));

shifter_right_tc #(.WIDTH(16), .SHIFT(16), .PAD_VALUE(1)) shifter_right_tc__width_16__shift_16__pad_1 (.start(start__shifter_right_tc__width_16__shift_16__pad_1));

shifter_right_tc #(.WIDTH(16), .SHIFT(17), .PAD_VALUE(1)) shifter_right_tc__width_16__shift_17__pad_1 (.start(start__shifter_right_tc__width_16__shift_17__pad_1));

shifter_right_tc #(.WIDTH(16), .SHIFT(24), .PAD_VALUE(1)) shifter_right_tc__width_16__shift_24__pad_1 (.start(start__shifter_right_tc__width_16__shift_24__pad_1));

shifter_right_tc #(.WIDTH(16), .SHIFT(31), .PAD_VALUE(1)) shifter_right_tc__width_16__shift_31__pad_1 (.start(start__shifter_right_tc__width_16__shift_31__pad_1));

shifter_right_tc #(.WIDTH(16), .SHIFT(32), .PAD_VALUE(1)) shifter_right_tc__width_16__shift_32__pad_1 (.start(start__shifter_right_tc__width_16__shift_32__pad_1));

shifter_right_tc #(.WIDTH(24), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_24__shift_0__pad_0 (.start(start__shifter_right_tc__width_24__shift_0__pad_0));

shifter_right_tc #(.WIDTH(24), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_24__shift_1__pad_0 (.start(start__shifter_right_tc__width_24__shift_1__pad_0));

shifter_right_tc #(.WIDTH(24), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_24__shift_2__pad_0 (.start(start__shifter_right_tc__width_24__shift_2__pad_0));

shifter_right_tc #(.WIDTH(24), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_24__shift_3__pad_0 (.start(start__shifter_right_tc__width_24__shift_3__pad_0));

shifter_right_tc #(.WIDTH(24), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_24__shift_4__pad_0 (.start(start__shifter_right_tc__width_24__shift_4__pad_0));

shifter_right_tc #(.WIDTH(24), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_24__shift_5__pad_0 (.start(start__shifter_right_tc__width_24__shift_5__pad_0));

shifter_right_tc #(.WIDTH(24), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_24__shift_6__pad_0 (.start(start__shifter_right_tc__width_24__shift_6__pad_0));

shifter_right_tc #(.WIDTH(24), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_24__shift_7__pad_0 (.start(start__shifter_right_tc__width_24__shift_7__pad_0));

shifter_right_tc #(.WIDTH(24), .SHIFT(12), .PAD_VALUE(0)) shifter_right_tc__width_24__shift_12__pad_0 (.start(start__shifter_right_tc__width_24__shift_12__pad_0));

shifter_right_tc #(.WIDTH(24), .SHIFT(23), .PAD_VALUE(0)) shifter_right_tc__width_24__shift_23__pad_0 (.start(start__shifter_right_tc__width_24__shift_23__pad_0));

shifter_right_tc #(.WIDTH(24), .SHIFT(24), .PAD_VALUE(0)) shifter_right_tc__width_24__shift_24__pad_0 (.start(start__shifter_right_tc__width_24__shift_24__pad_0));

shifter_right_tc #(.WIDTH(24), .SHIFT(25), .PAD_VALUE(0)) shifter_right_tc__width_24__shift_25__pad_0 (.start(start__shifter_right_tc__width_24__shift_25__pad_0));

shifter_right_tc #(.WIDTH(24), .SHIFT(36), .PAD_VALUE(0)) shifter_right_tc__width_24__shift_36__pad_0 (.start(start__shifter_right_tc__width_24__shift_36__pad_0));

shifter_right_tc #(.WIDTH(24), .SHIFT(47), .PAD_VALUE(0)) shifter_right_tc__width_24__shift_47__pad_0 (.start(start__shifter_right_tc__width_24__shift_47__pad_0));

shifter_right_tc #(.WIDTH(24), .SHIFT(48), .PAD_VALUE(0)) shifter_right_tc__width_24__shift_48__pad_0 (.start(start__shifter_right_tc__width_24__shift_48__pad_0));

shifter_right_tc #(.WIDTH(24), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_24__shift_0__pad_1 (.start(start__shifter_right_tc__width_24__shift_0__pad_1));

shifter_right_tc #(.WIDTH(24), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_24__shift_1__pad_1 (.start(start__shifter_right_tc__width_24__shift_1__pad_1));

shifter_right_tc #(.WIDTH(24), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_24__shift_2__pad_1 (.start(start__shifter_right_tc__width_24__shift_2__pad_1));

shifter_right_tc #(.WIDTH(24), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_24__shift_3__pad_1 (.start(start__shifter_right_tc__width_24__shift_3__pad_1));

shifter_right_tc #(.WIDTH(24), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_24__shift_4__pad_1 (.start(start__shifter_right_tc__width_24__shift_4__pad_1));

shifter_right_tc #(.WIDTH(24), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_24__shift_5__pad_1 (.start(start__shifter_right_tc__width_24__shift_5__pad_1));

shifter_right_tc #(.WIDTH(24), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_24__shift_6__pad_1 (.start(start__shifter_right_tc__width_24__shift_6__pad_1));

shifter_right_tc #(.WIDTH(24), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_24__shift_7__pad_1 (.start(start__shifter_right_tc__width_24__shift_7__pad_1));

shifter_right_tc #(.WIDTH(24), .SHIFT(12), .PAD_VALUE(1)) shifter_right_tc__width_24__shift_12__pad_1 (.start(start__shifter_right_tc__width_24__shift_12__pad_1));

shifter_right_tc #(.WIDTH(24), .SHIFT(23), .PAD_VALUE(1)) shifter_right_tc__width_24__shift_23__pad_1 (.start(start__shifter_right_tc__width_24__shift_23__pad_1));

shifter_right_tc #(.WIDTH(24), .SHIFT(24), .PAD_VALUE(1)) shifter_right_tc__width_24__shift_24__pad_1 (.start(start__shifter_right_tc__width_24__shift_24__pad_1));

shifter_right_tc #(.WIDTH(24), .SHIFT(25), .PAD_VALUE(1)) shifter_right_tc__width_24__shift_25__pad_1 (.start(start__shifter_right_tc__width_24__shift_25__pad_1));

shifter_right_tc #(.WIDTH(24), .SHIFT(36), .PAD_VALUE(1)) shifter_right_tc__width_24__shift_36__pad_1 (.start(start__shifter_right_tc__width_24__shift_36__pad_1));

shifter_right_tc #(.WIDTH(24), .SHIFT(47), .PAD_VALUE(1)) shifter_right_tc__width_24__shift_47__pad_1 (.start(start__shifter_right_tc__width_24__shift_47__pad_1));

shifter_right_tc #(.WIDTH(24), .SHIFT(48), .PAD_VALUE(1)) shifter_right_tc__width_24__shift_48__pad_1 (.start(start__shifter_right_tc__width_24__shift_48__pad_1));

shifter_right_tc #(.WIDTH(32), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_32__shift_0__pad_0 (.start(start__shifter_right_tc__width_32__shift_0__pad_0));

shifter_right_tc #(.WIDTH(32), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_32__shift_1__pad_0 (.start(start__shifter_right_tc__width_32__shift_1__pad_0));

shifter_right_tc #(.WIDTH(32), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_32__shift_2__pad_0 (.start(start__shifter_right_tc__width_32__shift_2__pad_0));

shifter_right_tc #(.WIDTH(32), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_32__shift_3__pad_0 (.start(start__shifter_right_tc__width_32__shift_3__pad_0));

shifter_right_tc #(.WIDTH(32), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_32__shift_4__pad_0 (.start(start__shifter_right_tc__width_32__shift_4__pad_0));

shifter_right_tc #(.WIDTH(32), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_32__shift_5__pad_0 (.start(start__shifter_right_tc__width_32__shift_5__pad_0));

shifter_right_tc #(.WIDTH(32), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_32__shift_6__pad_0 (.start(start__shifter_right_tc__width_32__shift_6__pad_0));

shifter_right_tc #(.WIDTH(32), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_32__shift_7__pad_0 (.start(start__shifter_right_tc__width_32__shift_7__pad_0));

shifter_right_tc #(.WIDTH(32), .SHIFT(16), .PAD_VALUE(0)) shifter_right_tc__width_32__shift_16__pad_0 (.start(start__shifter_right_tc__width_32__shift_16__pad_0));

shifter_right_tc #(.WIDTH(32), .SHIFT(31), .PAD_VALUE(0)) shifter_right_tc__width_32__shift_31__pad_0 (.start(start__shifter_right_tc__width_32__shift_31__pad_0));

shifter_right_tc #(.WIDTH(32), .SHIFT(32), .PAD_VALUE(0)) shifter_right_tc__width_32__shift_32__pad_0 (.start(start__shifter_right_tc__width_32__shift_32__pad_0));

shifter_right_tc #(.WIDTH(32), .SHIFT(33), .PAD_VALUE(0)) shifter_right_tc__width_32__shift_33__pad_0 (.start(start__shifter_right_tc__width_32__shift_33__pad_0));

shifter_right_tc #(.WIDTH(32), .SHIFT(48), .PAD_VALUE(0)) shifter_right_tc__width_32__shift_48__pad_0 (.start(start__shifter_right_tc__width_32__shift_48__pad_0));

shifter_right_tc #(.WIDTH(32), .SHIFT(63), .PAD_VALUE(0)) shifter_right_tc__width_32__shift_63__pad_0 (.start(start__shifter_right_tc__width_32__shift_63__pad_0));

shifter_right_tc #(.WIDTH(32), .SHIFT(64), .PAD_VALUE(0)) shifter_right_tc__width_32__shift_64__pad_0 (.start(start__shifter_right_tc__width_32__shift_64__pad_0));

shifter_right_tc #(.WIDTH(32), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_32__shift_0__pad_1 (.start(start__shifter_right_tc__width_32__shift_0__pad_1));

shifter_right_tc #(.WIDTH(32), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_32__shift_1__pad_1 (.start(start__shifter_right_tc__width_32__shift_1__pad_1));

shifter_right_tc #(.WIDTH(32), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_32__shift_2__pad_1 (.start(start__shifter_right_tc__width_32__shift_2__pad_1));

shifter_right_tc #(.WIDTH(32), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_32__shift_3__pad_1 (.start(start__shifter_right_tc__width_32__shift_3__pad_1));

shifter_right_tc #(.WIDTH(32), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_32__shift_4__pad_1 (.start(start__shifter_right_tc__width_32__shift_4__pad_1));

shifter_right_tc #(.WIDTH(32), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_32__shift_5__pad_1 (.start(start__shifter_right_tc__width_32__shift_5__pad_1));

shifter_right_tc #(.WIDTH(32), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_32__shift_6__pad_1 (.start(start__shifter_right_tc__width_32__shift_6__pad_1));

shifter_right_tc #(.WIDTH(32), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_32__shift_7__pad_1 (.start(start__shifter_right_tc__width_32__shift_7__pad_1));

shifter_right_tc #(.WIDTH(32), .SHIFT(16), .PAD_VALUE(1)) shifter_right_tc__width_32__shift_16__pad_1 (.start(start__shifter_right_tc__width_32__shift_16__pad_1));

shifter_right_tc #(.WIDTH(32), .SHIFT(31), .PAD_VALUE(1)) shifter_right_tc__width_32__shift_31__pad_1 (.start(start__shifter_right_tc__width_32__shift_31__pad_1));

shifter_right_tc #(.WIDTH(32), .SHIFT(32), .PAD_VALUE(1)) shifter_right_tc__width_32__shift_32__pad_1 (.start(start__shifter_right_tc__width_32__shift_32__pad_1));

shifter_right_tc #(.WIDTH(32), .SHIFT(33), .PAD_VALUE(1)) shifter_right_tc__width_32__shift_33__pad_1 (.start(start__shifter_right_tc__width_32__shift_33__pad_1));

shifter_right_tc #(.WIDTH(32), .SHIFT(48), .PAD_VALUE(1)) shifter_right_tc__width_32__shift_48__pad_1 (.start(start__shifter_right_tc__width_32__shift_48__pad_1));

shifter_right_tc #(.WIDTH(32), .SHIFT(63), .PAD_VALUE(1)) shifter_right_tc__width_32__shift_63__pad_1 (.start(start__shifter_right_tc__width_32__shift_63__pad_1));

shifter_right_tc #(.WIDTH(32), .SHIFT(64), .PAD_VALUE(1)) shifter_right_tc__width_32__shift_64__pad_1 (.start(start__shifter_right_tc__width_32__shift_64__pad_1));

shifter_right_tc #(.WIDTH(48), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_48__shift_0__pad_0 (.start(start__shifter_right_tc__width_48__shift_0__pad_0));

shifter_right_tc #(.WIDTH(48), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_48__shift_1__pad_0 (.start(start__shifter_right_tc__width_48__shift_1__pad_0));

shifter_right_tc #(.WIDTH(48), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_48__shift_2__pad_0 (.start(start__shifter_right_tc__width_48__shift_2__pad_0));

shifter_right_tc #(.WIDTH(48), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_48__shift_3__pad_0 (.start(start__shifter_right_tc__width_48__shift_3__pad_0));

shifter_right_tc #(.WIDTH(48), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_48__shift_4__pad_0 (.start(start__shifter_right_tc__width_48__shift_4__pad_0));

shifter_right_tc #(.WIDTH(48), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_48__shift_5__pad_0 (.start(start__shifter_right_tc__width_48__shift_5__pad_0));

shifter_right_tc #(.WIDTH(48), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_48__shift_6__pad_0 (.start(start__shifter_right_tc__width_48__shift_6__pad_0));

shifter_right_tc #(.WIDTH(48), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_48__shift_7__pad_0 (.start(start__shifter_right_tc__width_48__shift_7__pad_0));

shifter_right_tc #(.WIDTH(48), .SHIFT(24), .PAD_VALUE(0)) shifter_right_tc__width_48__shift_24__pad_0 (.start(start__shifter_right_tc__width_48__shift_24__pad_0));

shifter_right_tc #(.WIDTH(48), .SHIFT(47), .PAD_VALUE(0)) shifter_right_tc__width_48__shift_47__pad_0 (.start(start__shifter_right_tc__width_48__shift_47__pad_0));

shifter_right_tc #(.WIDTH(48), .SHIFT(48), .PAD_VALUE(0)) shifter_right_tc__width_48__shift_48__pad_0 (.start(start__shifter_right_tc__width_48__shift_48__pad_0));

shifter_right_tc #(.WIDTH(48), .SHIFT(49), .PAD_VALUE(0)) shifter_right_tc__width_48__shift_49__pad_0 (.start(start__shifter_right_tc__width_48__shift_49__pad_0));

shifter_right_tc #(.WIDTH(48), .SHIFT(72), .PAD_VALUE(0)) shifter_right_tc__width_48__shift_72__pad_0 (.start(start__shifter_right_tc__width_48__shift_72__pad_0));

shifter_right_tc #(.WIDTH(48), .SHIFT(95), .PAD_VALUE(0)) shifter_right_tc__width_48__shift_95__pad_0 (.start(start__shifter_right_tc__width_48__shift_95__pad_0));

shifter_right_tc #(.WIDTH(48), .SHIFT(96), .PAD_VALUE(0)) shifter_right_tc__width_48__shift_96__pad_0 (.start(start__shifter_right_tc__width_48__shift_96__pad_0));

shifter_right_tc #(.WIDTH(48), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_48__shift_0__pad_1 (.start(start__shifter_right_tc__width_48__shift_0__pad_1));

shifter_right_tc #(.WIDTH(48), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_48__shift_1__pad_1 (.start(start__shifter_right_tc__width_48__shift_1__pad_1));

shifter_right_tc #(.WIDTH(48), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_48__shift_2__pad_1 (.start(start__shifter_right_tc__width_48__shift_2__pad_1));

shifter_right_tc #(.WIDTH(48), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_48__shift_3__pad_1 (.start(start__shifter_right_tc__width_48__shift_3__pad_1));

shifter_right_tc #(.WIDTH(48), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_48__shift_4__pad_1 (.start(start__shifter_right_tc__width_48__shift_4__pad_1));

shifter_right_tc #(.WIDTH(48), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_48__shift_5__pad_1 (.start(start__shifter_right_tc__width_48__shift_5__pad_1));

shifter_right_tc #(.WIDTH(48), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_48__shift_6__pad_1 (.start(start__shifter_right_tc__width_48__shift_6__pad_1));

shifter_right_tc #(.WIDTH(48), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_48__shift_7__pad_1 (.start(start__shifter_right_tc__width_48__shift_7__pad_1));

shifter_right_tc #(.WIDTH(48), .SHIFT(24), .PAD_VALUE(1)) shifter_right_tc__width_48__shift_24__pad_1 (.start(start__shifter_right_tc__width_48__shift_24__pad_1));

shifter_right_tc #(.WIDTH(48), .SHIFT(47), .PAD_VALUE(1)) shifter_right_tc__width_48__shift_47__pad_1 (.start(start__shifter_right_tc__width_48__shift_47__pad_1));

shifter_right_tc #(.WIDTH(48), .SHIFT(48), .PAD_VALUE(1)) shifter_right_tc__width_48__shift_48__pad_1 (.start(start__shifter_right_tc__width_48__shift_48__pad_1));

shifter_right_tc #(.WIDTH(48), .SHIFT(49), .PAD_VALUE(1)) shifter_right_tc__width_48__shift_49__pad_1 (.start(start__shifter_right_tc__width_48__shift_49__pad_1));

shifter_right_tc #(.WIDTH(48), .SHIFT(72), .PAD_VALUE(1)) shifter_right_tc__width_48__shift_72__pad_1 (.start(start__shifter_right_tc__width_48__shift_72__pad_1));

shifter_right_tc #(.WIDTH(48), .SHIFT(95), .PAD_VALUE(1)) shifter_right_tc__width_48__shift_95__pad_1 (.start(start__shifter_right_tc__width_48__shift_95__pad_1));

shifter_right_tc #(.WIDTH(48), .SHIFT(96), .PAD_VALUE(1)) shifter_right_tc__width_48__shift_96__pad_1 (.start(start__shifter_right_tc__width_48__shift_96__pad_1));

shifter_right_tc #(.WIDTH(64), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_64__shift_0__pad_0 (.start(start__shifter_right_tc__width_64__shift_0__pad_0));

shifter_right_tc #(.WIDTH(64), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_64__shift_1__pad_0 (.start(start__shifter_right_tc__width_64__shift_1__pad_0));

shifter_right_tc #(.WIDTH(64), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_64__shift_2__pad_0 (.start(start__shifter_right_tc__width_64__shift_2__pad_0));

shifter_right_tc #(.WIDTH(64), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_64__shift_3__pad_0 (.start(start__shifter_right_tc__width_64__shift_3__pad_0));

shifter_right_tc #(.WIDTH(64), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_64__shift_4__pad_0 (.start(start__shifter_right_tc__width_64__shift_4__pad_0));

shifter_right_tc #(.WIDTH(64), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_64__shift_5__pad_0 (.start(start__shifter_right_tc__width_64__shift_5__pad_0));

shifter_right_tc #(.WIDTH(64), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_64__shift_6__pad_0 (.start(start__shifter_right_tc__width_64__shift_6__pad_0));

shifter_right_tc #(.WIDTH(64), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_64__shift_7__pad_0 (.start(start__shifter_right_tc__width_64__shift_7__pad_0));

shifter_right_tc #(.WIDTH(64), .SHIFT(32), .PAD_VALUE(0)) shifter_right_tc__width_64__shift_32__pad_0 (.start(start__shifter_right_tc__width_64__shift_32__pad_0));

shifter_right_tc #(.WIDTH(64), .SHIFT(63), .PAD_VALUE(0)) shifter_right_tc__width_64__shift_63__pad_0 (.start(start__shifter_right_tc__width_64__shift_63__pad_0));

shifter_right_tc #(.WIDTH(64), .SHIFT(64), .PAD_VALUE(0)) shifter_right_tc__width_64__shift_64__pad_0 (.start(start__shifter_right_tc__width_64__shift_64__pad_0));

shifter_right_tc #(.WIDTH(64), .SHIFT(65), .PAD_VALUE(0)) shifter_right_tc__width_64__shift_65__pad_0 (.start(start__shifter_right_tc__width_64__shift_65__pad_0));

shifter_right_tc #(.WIDTH(64), .SHIFT(96), .PAD_VALUE(0)) shifter_right_tc__width_64__shift_96__pad_0 (.start(start__shifter_right_tc__width_64__shift_96__pad_0));

shifter_right_tc #(.WIDTH(64), .SHIFT(127), .PAD_VALUE(0)) shifter_right_tc__width_64__shift_127__pad_0 (.start(start__shifter_right_tc__width_64__shift_127__pad_0));

shifter_right_tc #(.WIDTH(64), .SHIFT(128), .PAD_VALUE(0)) shifter_right_tc__width_64__shift_128__pad_0 (.start(start__shifter_right_tc__width_64__shift_128__pad_0));

shifter_right_tc #(.WIDTH(64), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_64__shift_0__pad_1 (.start(start__shifter_right_tc__width_64__shift_0__pad_1));

shifter_right_tc #(.WIDTH(64), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_64__shift_1__pad_1 (.start(start__shifter_right_tc__width_64__shift_1__pad_1));

shifter_right_tc #(.WIDTH(64), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_64__shift_2__pad_1 (.start(start__shifter_right_tc__width_64__shift_2__pad_1));

shifter_right_tc #(.WIDTH(64), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_64__shift_3__pad_1 (.start(start__shifter_right_tc__width_64__shift_3__pad_1));

shifter_right_tc #(.WIDTH(64), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_64__shift_4__pad_1 (.start(start__shifter_right_tc__width_64__shift_4__pad_1));

shifter_right_tc #(.WIDTH(64), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_64__shift_5__pad_1 (.start(start__shifter_right_tc__width_64__shift_5__pad_1));

shifter_right_tc #(.WIDTH(64), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_64__shift_6__pad_1 (.start(start__shifter_right_tc__width_64__shift_6__pad_1));

shifter_right_tc #(.WIDTH(64), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_64__shift_7__pad_1 (.start(start__shifter_right_tc__width_64__shift_7__pad_1));

shifter_right_tc #(.WIDTH(64), .SHIFT(32), .PAD_VALUE(1)) shifter_right_tc__width_64__shift_32__pad_1 (.start(start__shifter_right_tc__width_64__shift_32__pad_1));

shifter_right_tc #(.WIDTH(64), .SHIFT(63), .PAD_VALUE(1)) shifter_right_tc__width_64__shift_63__pad_1 (.start(start__shifter_right_tc__width_64__shift_63__pad_1));

shifter_right_tc #(.WIDTH(64), .SHIFT(64), .PAD_VALUE(1)) shifter_right_tc__width_64__shift_64__pad_1 (.start(start__shifter_right_tc__width_64__shift_64__pad_1));

shifter_right_tc #(.WIDTH(64), .SHIFT(65), .PAD_VALUE(1)) shifter_right_tc__width_64__shift_65__pad_1 (.start(start__shifter_right_tc__width_64__shift_65__pad_1));

shifter_right_tc #(.WIDTH(64), .SHIFT(96), .PAD_VALUE(1)) shifter_right_tc__width_64__shift_96__pad_1 (.start(start__shifter_right_tc__width_64__shift_96__pad_1));

shifter_right_tc #(.WIDTH(64), .SHIFT(127), .PAD_VALUE(1)) shifter_right_tc__width_64__shift_127__pad_1 (.start(start__shifter_right_tc__width_64__shift_127__pad_1));

shifter_right_tc #(.WIDTH(64), .SHIFT(128), .PAD_VALUE(1)) shifter_right_tc__width_64__shift_128__pad_1 (.start(start__shifter_right_tc__width_64__shift_128__pad_1));

shifter_right_tc #(.WIDTH(128), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_128__shift_0__pad_0 (.start(start__shifter_right_tc__width_128__shift_0__pad_0));

shifter_right_tc #(.WIDTH(128), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_128__shift_1__pad_0 (.start(start__shifter_right_tc__width_128__shift_1__pad_0));

shifter_right_tc #(.WIDTH(128), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_128__shift_2__pad_0 (.start(start__shifter_right_tc__width_128__shift_2__pad_0));

shifter_right_tc #(.WIDTH(128), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_128__shift_3__pad_0 (.start(start__shifter_right_tc__width_128__shift_3__pad_0));

shifter_right_tc #(.WIDTH(128), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_128__shift_4__pad_0 (.start(start__shifter_right_tc__width_128__shift_4__pad_0));

shifter_right_tc #(.WIDTH(128), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_128__shift_5__pad_0 (.start(start__shifter_right_tc__width_128__shift_5__pad_0));

shifter_right_tc #(.WIDTH(128), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_128__shift_6__pad_0 (.start(start__shifter_right_tc__width_128__shift_6__pad_0));

shifter_right_tc #(.WIDTH(128), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_128__shift_7__pad_0 (.start(start__shifter_right_tc__width_128__shift_7__pad_0));

shifter_right_tc #(.WIDTH(128), .SHIFT(64), .PAD_VALUE(0)) shifter_right_tc__width_128__shift_64__pad_0 (.start(start__shifter_right_tc__width_128__shift_64__pad_0));

shifter_right_tc #(.WIDTH(128), .SHIFT(127), .PAD_VALUE(0)) shifter_right_tc__width_128__shift_127__pad_0 (.start(start__shifter_right_tc__width_128__shift_127__pad_0));

shifter_right_tc #(.WIDTH(128), .SHIFT(128), .PAD_VALUE(0)) shifter_right_tc__width_128__shift_128__pad_0 (.start(start__shifter_right_tc__width_128__shift_128__pad_0));

shifter_right_tc #(.WIDTH(128), .SHIFT(129), .PAD_VALUE(0)) shifter_right_tc__width_128__shift_129__pad_0 (.start(start__shifter_right_tc__width_128__shift_129__pad_0));

shifter_right_tc #(.WIDTH(128), .SHIFT(192), .PAD_VALUE(0)) shifter_right_tc__width_128__shift_192__pad_0 (.start(start__shifter_right_tc__width_128__shift_192__pad_0));

shifter_right_tc #(.WIDTH(128), .SHIFT(255), .PAD_VALUE(0)) shifter_right_tc__width_128__shift_255__pad_0 (.start(start__shifter_right_tc__width_128__shift_255__pad_0));

shifter_right_tc #(.WIDTH(128), .SHIFT(256), .PAD_VALUE(0)) shifter_right_tc__width_128__shift_256__pad_0 (.start(start__shifter_right_tc__width_128__shift_256__pad_0));

shifter_right_tc #(.WIDTH(128), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_128__shift_0__pad_1 (.start(start__shifter_right_tc__width_128__shift_0__pad_1));

shifter_right_tc #(.WIDTH(128), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_128__shift_1__pad_1 (.start(start__shifter_right_tc__width_128__shift_1__pad_1));

shifter_right_tc #(.WIDTH(128), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_128__shift_2__pad_1 (.start(start__shifter_right_tc__width_128__shift_2__pad_1));

shifter_right_tc #(.WIDTH(128), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_128__shift_3__pad_1 (.start(start__shifter_right_tc__width_128__shift_3__pad_1));

shifter_right_tc #(.WIDTH(128), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_128__shift_4__pad_1 (.start(start__shifter_right_tc__width_128__shift_4__pad_1));

shifter_right_tc #(.WIDTH(128), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_128__shift_5__pad_1 (.start(start__shifter_right_tc__width_128__shift_5__pad_1));

shifter_right_tc #(.WIDTH(128), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_128__shift_6__pad_1 (.start(start__shifter_right_tc__width_128__shift_6__pad_1));

shifter_right_tc #(.WIDTH(128), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_128__shift_7__pad_1 (.start(start__shifter_right_tc__width_128__shift_7__pad_1));

shifter_right_tc #(.WIDTH(128), .SHIFT(64), .PAD_VALUE(1)) shifter_right_tc__width_128__shift_64__pad_1 (.start(start__shifter_right_tc__width_128__shift_64__pad_1));

shifter_right_tc #(.WIDTH(128), .SHIFT(127), .PAD_VALUE(1)) shifter_right_tc__width_128__shift_127__pad_1 (.start(start__shifter_right_tc__width_128__shift_127__pad_1));

shifter_right_tc #(.WIDTH(128), .SHIFT(128), .PAD_VALUE(1)) shifter_right_tc__width_128__shift_128__pad_1 (.start(start__shifter_right_tc__width_128__shift_128__pad_1));

shifter_right_tc #(.WIDTH(128), .SHIFT(129), .PAD_VALUE(1)) shifter_right_tc__width_128__shift_129__pad_1 (.start(start__shifter_right_tc__width_128__shift_129__pad_1));

shifter_right_tc #(.WIDTH(128), .SHIFT(192), .PAD_VALUE(1)) shifter_right_tc__width_128__shift_192__pad_1 (.start(start__shifter_right_tc__width_128__shift_192__pad_1));

shifter_right_tc #(.WIDTH(128), .SHIFT(255), .PAD_VALUE(1)) shifter_right_tc__width_128__shift_255__pad_1 (.start(start__shifter_right_tc__width_128__shift_255__pad_1));

shifter_right_tc #(.WIDTH(128), .SHIFT(256), .PAD_VALUE(1)) shifter_right_tc__width_128__shift_256__pad_1 (.start(start__shifter_right_tc__width_128__shift_256__pad_1));

shifter_right_tc #(.WIDTH(256), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_256__shift_0__pad_0 (.start(start__shifter_right_tc__width_256__shift_0__pad_0));

shifter_right_tc #(.WIDTH(256), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_256__shift_1__pad_0 (.start(start__shifter_right_tc__width_256__shift_1__pad_0));

shifter_right_tc #(.WIDTH(256), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_256__shift_2__pad_0 (.start(start__shifter_right_tc__width_256__shift_2__pad_0));

shifter_right_tc #(.WIDTH(256), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_256__shift_3__pad_0 (.start(start__shifter_right_tc__width_256__shift_3__pad_0));

shifter_right_tc #(.WIDTH(256), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_256__shift_4__pad_0 (.start(start__shifter_right_tc__width_256__shift_4__pad_0));

shifter_right_tc #(.WIDTH(256), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_256__shift_5__pad_0 (.start(start__shifter_right_tc__width_256__shift_5__pad_0));

shifter_right_tc #(.WIDTH(256), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_256__shift_6__pad_0 (.start(start__shifter_right_tc__width_256__shift_6__pad_0));

shifter_right_tc #(.WIDTH(256), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_256__shift_7__pad_0 (.start(start__shifter_right_tc__width_256__shift_7__pad_0));

shifter_right_tc #(.WIDTH(256), .SHIFT(128), .PAD_VALUE(0)) shifter_right_tc__width_256__shift_128__pad_0 (.start(start__shifter_right_tc__width_256__shift_128__pad_0));

shifter_right_tc #(.WIDTH(256), .SHIFT(255), .PAD_VALUE(0)) shifter_right_tc__width_256__shift_255__pad_0 (.start(start__shifter_right_tc__width_256__shift_255__pad_0));

shifter_right_tc #(.WIDTH(256), .SHIFT(256), .PAD_VALUE(0)) shifter_right_tc__width_256__shift_256__pad_0 (.start(start__shifter_right_tc__width_256__shift_256__pad_0));

shifter_right_tc #(.WIDTH(256), .SHIFT(257), .PAD_VALUE(0)) shifter_right_tc__width_256__shift_257__pad_0 (.start(start__shifter_right_tc__width_256__shift_257__pad_0));

shifter_right_tc #(.WIDTH(256), .SHIFT(384), .PAD_VALUE(0)) shifter_right_tc__width_256__shift_384__pad_0 (.start(start__shifter_right_tc__width_256__shift_384__pad_0));

shifter_right_tc #(.WIDTH(256), .SHIFT(511), .PAD_VALUE(0)) shifter_right_tc__width_256__shift_511__pad_0 (.start(start__shifter_right_tc__width_256__shift_511__pad_0));

shifter_right_tc #(.WIDTH(256), .SHIFT(512), .PAD_VALUE(0)) shifter_right_tc__width_256__shift_512__pad_0 (.start(start__shifter_right_tc__width_256__shift_512__pad_0));

shifter_right_tc #(.WIDTH(256), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_256__shift_0__pad_1 (.start(start__shifter_right_tc__width_256__shift_0__pad_1));

shifter_right_tc #(.WIDTH(256), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_256__shift_1__pad_1 (.start(start__shifter_right_tc__width_256__shift_1__pad_1));

shifter_right_tc #(.WIDTH(256), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_256__shift_2__pad_1 (.start(start__shifter_right_tc__width_256__shift_2__pad_1));

shifter_right_tc #(.WIDTH(256), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_256__shift_3__pad_1 (.start(start__shifter_right_tc__width_256__shift_3__pad_1));

shifter_right_tc #(.WIDTH(256), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_256__shift_4__pad_1 (.start(start__shifter_right_tc__width_256__shift_4__pad_1));

shifter_right_tc #(.WIDTH(256), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_256__shift_5__pad_1 (.start(start__shifter_right_tc__width_256__shift_5__pad_1));

shifter_right_tc #(.WIDTH(256), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_256__shift_6__pad_1 (.start(start__shifter_right_tc__width_256__shift_6__pad_1));

shifter_right_tc #(.WIDTH(256), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_256__shift_7__pad_1 (.start(start__shifter_right_tc__width_256__shift_7__pad_1));

shifter_right_tc #(.WIDTH(256), .SHIFT(128), .PAD_VALUE(1)) shifter_right_tc__width_256__shift_128__pad_1 (.start(start__shifter_right_tc__width_256__shift_128__pad_1));

shifter_right_tc #(.WIDTH(256), .SHIFT(255), .PAD_VALUE(1)) shifter_right_tc__width_256__shift_255__pad_1 (.start(start__shifter_right_tc__width_256__shift_255__pad_1));

shifter_right_tc #(.WIDTH(256), .SHIFT(256), .PAD_VALUE(1)) shifter_right_tc__width_256__shift_256__pad_1 (.start(start__shifter_right_tc__width_256__shift_256__pad_1));

shifter_right_tc #(.WIDTH(256), .SHIFT(257), .PAD_VALUE(1)) shifter_right_tc__width_256__shift_257__pad_1 (.start(start__shifter_right_tc__width_256__shift_257__pad_1));

shifter_right_tc #(.WIDTH(256), .SHIFT(384), .PAD_VALUE(1)) shifter_right_tc__width_256__shift_384__pad_1 (.start(start__shifter_right_tc__width_256__shift_384__pad_1));

shifter_right_tc #(.WIDTH(256), .SHIFT(511), .PAD_VALUE(1)) shifter_right_tc__width_256__shift_511__pad_1 (.start(start__shifter_right_tc__width_256__shift_511__pad_1));

shifter_right_tc #(.WIDTH(256), .SHIFT(512), .PAD_VALUE(1)) shifter_right_tc__width_256__shift_512__pad_1 (.start(start__shifter_right_tc__width_256__shift_512__pad_1));

shifter_right_tc #(.WIDTH(512), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_512__shift_0__pad_0 (.start(start__shifter_right_tc__width_512__shift_0__pad_0));

shifter_right_tc #(.WIDTH(512), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_512__shift_1__pad_0 (.start(start__shifter_right_tc__width_512__shift_1__pad_0));

shifter_right_tc #(.WIDTH(512), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_512__shift_2__pad_0 (.start(start__shifter_right_tc__width_512__shift_2__pad_0));

shifter_right_tc #(.WIDTH(512), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_512__shift_3__pad_0 (.start(start__shifter_right_tc__width_512__shift_3__pad_0));

shifter_right_tc #(.WIDTH(512), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_512__shift_4__pad_0 (.start(start__shifter_right_tc__width_512__shift_4__pad_0));

shifter_right_tc #(.WIDTH(512), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_512__shift_5__pad_0 (.start(start__shifter_right_tc__width_512__shift_5__pad_0));

shifter_right_tc #(.WIDTH(512), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_512__shift_6__pad_0 (.start(start__shifter_right_tc__width_512__shift_6__pad_0));

shifter_right_tc #(.WIDTH(512), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_512__shift_7__pad_0 (.start(start__shifter_right_tc__width_512__shift_7__pad_0));

shifter_right_tc #(.WIDTH(512), .SHIFT(256), .PAD_VALUE(0)) shifter_right_tc__width_512__shift_256__pad_0 (.start(start__shifter_right_tc__width_512__shift_256__pad_0));

shifter_right_tc #(.WIDTH(512), .SHIFT(511), .PAD_VALUE(0)) shifter_right_tc__width_512__shift_511__pad_0 (.start(start__shifter_right_tc__width_512__shift_511__pad_0));

shifter_right_tc #(.WIDTH(512), .SHIFT(512), .PAD_VALUE(0)) shifter_right_tc__width_512__shift_512__pad_0 (.start(start__shifter_right_tc__width_512__shift_512__pad_0));

shifter_right_tc #(.WIDTH(512), .SHIFT(513), .PAD_VALUE(0)) shifter_right_tc__width_512__shift_513__pad_0 (.start(start__shifter_right_tc__width_512__shift_513__pad_0));

shifter_right_tc #(.WIDTH(512), .SHIFT(768), .PAD_VALUE(0)) shifter_right_tc__width_512__shift_768__pad_0 (.start(start__shifter_right_tc__width_512__shift_768__pad_0));

shifter_right_tc #(.WIDTH(512), .SHIFT(1023), .PAD_VALUE(0)) shifter_right_tc__width_512__shift_1023__pad_0 (.start(start__shifter_right_tc__width_512__shift_1023__pad_0));

shifter_right_tc #(.WIDTH(512), .SHIFT(1024), .PAD_VALUE(0)) shifter_right_tc__width_512__shift_1024__pad_0 (.start(start__shifter_right_tc__width_512__shift_1024__pad_0));

shifter_right_tc #(.WIDTH(512), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_512__shift_0__pad_1 (.start(start__shifter_right_tc__width_512__shift_0__pad_1));

shifter_right_tc #(.WIDTH(512), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_512__shift_1__pad_1 (.start(start__shifter_right_tc__width_512__shift_1__pad_1));

shifter_right_tc #(.WIDTH(512), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_512__shift_2__pad_1 (.start(start__shifter_right_tc__width_512__shift_2__pad_1));

shifter_right_tc #(.WIDTH(512), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_512__shift_3__pad_1 (.start(start__shifter_right_tc__width_512__shift_3__pad_1));

shifter_right_tc #(.WIDTH(512), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_512__shift_4__pad_1 (.start(start__shifter_right_tc__width_512__shift_4__pad_1));

shifter_right_tc #(.WIDTH(512), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_512__shift_5__pad_1 (.start(start__shifter_right_tc__width_512__shift_5__pad_1));

shifter_right_tc #(.WIDTH(512), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_512__shift_6__pad_1 (.start(start__shifter_right_tc__width_512__shift_6__pad_1));

shifter_right_tc #(.WIDTH(512), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_512__shift_7__pad_1 (.start(start__shifter_right_tc__width_512__shift_7__pad_1));

shifter_right_tc #(.WIDTH(512), .SHIFT(256), .PAD_VALUE(1)) shifter_right_tc__width_512__shift_256__pad_1 (.start(start__shifter_right_tc__width_512__shift_256__pad_1));

shifter_right_tc #(.WIDTH(512), .SHIFT(511), .PAD_VALUE(1)) shifter_right_tc__width_512__shift_511__pad_1 (.start(start__shifter_right_tc__width_512__shift_511__pad_1));

shifter_right_tc #(.WIDTH(512), .SHIFT(512), .PAD_VALUE(1)) shifter_right_tc__width_512__shift_512__pad_1 (.start(start__shifter_right_tc__width_512__shift_512__pad_1));

shifter_right_tc #(.WIDTH(512), .SHIFT(513), .PAD_VALUE(1)) shifter_right_tc__width_512__shift_513__pad_1 (.start(start__shifter_right_tc__width_512__shift_513__pad_1));

shifter_right_tc #(.WIDTH(512), .SHIFT(768), .PAD_VALUE(1)) shifter_right_tc__width_512__shift_768__pad_1 (.start(start__shifter_right_tc__width_512__shift_768__pad_1));

shifter_right_tc #(.WIDTH(512), .SHIFT(1023), .PAD_VALUE(1)) shifter_right_tc__width_512__shift_1023__pad_1 (.start(start__shifter_right_tc__width_512__shift_1023__pad_1));

shifter_right_tc #(.WIDTH(512), .SHIFT(1024), .PAD_VALUE(1)) shifter_right_tc__width_512__shift_1024__pad_1 (.start(start__shifter_right_tc__width_512__shift_1024__pad_1));

shifter_right_tc #(.WIDTH(1024), .SHIFT(0), .PAD_VALUE(0)) shifter_right_tc__width_1024__shift_0__pad_0 (.start(start__shifter_right_tc__width_1024__shift_0__pad_0));

shifter_right_tc #(.WIDTH(1024), .SHIFT(1), .PAD_VALUE(0)) shifter_right_tc__width_1024__shift_1__pad_0 (.start(start__shifter_right_tc__width_1024__shift_1__pad_0));

shifter_right_tc #(.WIDTH(1024), .SHIFT(2), .PAD_VALUE(0)) shifter_right_tc__width_1024__shift_2__pad_0 (.start(start__shifter_right_tc__width_1024__shift_2__pad_0));

shifter_right_tc #(.WIDTH(1024), .SHIFT(3), .PAD_VALUE(0)) shifter_right_tc__width_1024__shift_3__pad_0 (.start(start__shifter_right_tc__width_1024__shift_3__pad_0));

shifter_right_tc #(.WIDTH(1024), .SHIFT(4), .PAD_VALUE(0)) shifter_right_tc__width_1024__shift_4__pad_0 (.start(start__shifter_right_tc__width_1024__shift_4__pad_0));

shifter_right_tc #(.WIDTH(1024), .SHIFT(5), .PAD_VALUE(0)) shifter_right_tc__width_1024__shift_5__pad_0 (.start(start__shifter_right_tc__width_1024__shift_5__pad_0));

shifter_right_tc #(.WIDTH(1024), .SHIFT(6), .PAD_VALUE(0)) shifter_right_tc__width_1024__shift_6__pad_0 (.start(start__shifter_right_tc__width_1024__shift_6__pad_0));

shifter_right_tc #(.WIDTH(1024), .SHIFT(7), .PAD_VALUE(0)) shifter_right_tc__width_1024__shift_7__pad_0 (.start(start__shifter_right_tc__width_1024__shift_7__pad_0));

shifter_right_tc #(.WIDTH(1024), .SHIFT(512), .PAD_VALUE(0)) shifter_right_tc__width_1024__shift_512__pad_0 (.start(start__shifter_right_tc__width_1024__shift_512__pad_0));

shifter_right_tc #(.WIDTH(1024), .SHIFT(1023), .PAD_VALUE(0)) shifter_right_tc__width_1024__shift_1023__pad_0 (.start(start__shifter_right_tc__width_1024__shift_1023__pad_0));

shifter_right_tc #(.WIDTH(1024), .SHIFT(1024), .PAD_VALUE(0)) shifter_right_tc__width_1024__shift_1024__pad_0 (.start(start__shifter_right_tc__width_1024__shift_1024__pad_0));

shifter_right_tc #(.WIDTH(1024), .SHIFT(1025), .PAD_VALUE(0)) shifter_right_tc__width_1024__shift_1025__pad_0 (.start(start__shifter_right_tc__width_1024__shift_1025__pad_0));

shifter_right_tc #(.WIDTH(1024), .SHIFT(1536), .PAD_VALUE(0)) shifter_right_tc__width_1024__shift_1536__pad_0 (.start(start__shifter_right_tc__width_1024__shift_1536__pad_0));

shifter_right_tc #(.WIDTH(1024), .SHIFT(2047), .PAD_VALUE(0)) shifter_right_tc__width_1024__shift_2047__pad_0 (.start(start__shifter_right_tc__width_1024__shift_2047__pad_0));

shifter_right_tc #(.WIDTH(1024), .SHIFT(2048), .PAD_VALUE(0)) shifter_right_tc__width_1024__shift_2048__pad_0 (.start(start__shifter_right_tc__width_1024__shift_2048__pad_0));

shifter_right_tc #(.WIDTH(1024), .SHIFT(0), .PAD_VALUE(1)) shifter_right_tc__width_1024__shift_0__pad_1 (.start(start__shifter_right_tc__width_1024__shift_0__pad_1));

shifter_right_tc #(.WIDTH(1024), .SHIFT(1), .PAD_VALUE(1)) shifter_right_tc__width_1024__shift_1__pad_1 (.start(start__shifter_right_tc__width_1024__shift_1__pad_1));

shifter_right_tc #(.WIDTH(1024), .SHIFT(2), .PAD_VALUE(1)) shifter_right_tc__width_1024__shift_2__pad_1 (.start(start__shifter_right_tc__width_1024__shift_2__pad_1));

shifter_right_tc #(.WIDTH(1024), .SHIFT(3), .PAD_VALUE(1)) shifter_right_tc__width_1024__shift_3__pad_1 (.start(start__shifter_right_tc__width_1024__shift_3__pad_1));

shifter_right_tc #(.WIDTH(1024), .SHIFT(4), .PAD_VALUE(1)) shifter_right_tc__width_1024__shift_4__pad_1 (.start(start__shifter_right_tc__width_1024__shift_4__pad_1));

shifter_right_tc #(.WIDTH(1024), .SHIFT(5), .PAD_VALUE(1)) shifter_right_tc__width_1024__shift_5__pad_1 (.start(start__shifter_right_tc__width_1024__shift_5__pad_1));

shifter_right_tc #(.WIDTH(1024), .SHIFT(6), .PAD_VALUE(1)) shifter_right_tc__width_1024__shift_6__pad_1 (.start(start__shifter_right_tc__width_1024__shift_6__pad_1));

shifter_right_tc #(.WIDTH(1024), .SHIFT(7), .PAD_VALUE(1)) shifter_right_tc__width_1024__shift_7__pad_1 (.start(start__shifter_right_tc__width_1024__shift_7__pad_1));

shifter_right_tc #(.WIDTH(1024), .SHIFT(512), .PAD_VALUE(1)) shifter_right_tc__width_1024__shift_512__pad_1 (.start(start__shifter_right_tc__width_1024__shift_512__pad_1));

shifter_right_tc #(.WIDTH(1024), .SHIFT(1023), .PAD_VALUE(1)) shifter_right_tc__width_1024__shift_1023__pad_1 (.start(start__shifter_right_tc__width_1024__shift_1023__pad_1));

shifter_right_tc #(.WIDTH(1024), .SHIFT(1024), .PAD_VALUE(1)) shifter_right_tc__width_1024__shift_1024__pad_1 (.start(start__shifter_right_tc__width_1024__shift_1024__pad_1));

shifter_right_tc #(.WIDTH(1024), .SHIFT(1025), .PAD_VALUE(1)) shifter_right_tc__width_1024__shift_1025__pad_1 (.start(start__shifter_right_tc__width_1024__shift_1025__pad_1));

shifter_right_tc #(.WIDTH(1024), .SHIFT(1536), .PAD_VALUE(1)) shifter_right_tc__width_1024__shift_1536__pad_1 (.start(start__shifter_right_tc__width_1024__shift_1536__pad_1));

shifter_right_tc #(.WIDTH(1024), .SHIFT(2047), .PAD_VALUE(1)) shifter_right_tc__width_1024__shift_2047__pad_1 (.start(start__shifter_right_tc__width_1024__shift_2047__pad_1));

shifter_right_tc #(.WIDTH(1024), .SHIFT(2048), .PAD_VALUE(1)) shifter_right_tc__width_1024__shift_2048__pad_1 (.start(start__shifter_right_tc__width_1024__shift_2048__pad_1));


initial begin
  // Log waves
  $dumpfile("shifter_right.tb.vcd");


  $dumpvars(0,shifter_right_tc__width_1__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_1__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_1__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_1__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_2__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_2__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_2__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_2__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_2__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_2__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_2__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_2__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_3__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_3__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_3__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_3__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_3__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_3__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_3__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_3__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_3__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_3__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_3__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_3__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_4__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_4__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_4__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_4__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_4__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_4__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_4__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_4__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_4__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_4__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_4__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_4__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_4__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_4__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_4__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_4__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_5__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_5__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_5__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_5__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_5__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_5__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_5__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_5__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_5__shift_8__pad_0);

  $dumpvars(0,shifter_right_tc__width_5__shift_9__pad_0);

  $dumpvars(0,shifter_right_tc__width_5__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_5__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_5__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_5__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_5__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_5__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_5__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_5__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_5__shift_8__pad_1);

  $dumpvars(0,shifter_right_tc__width_5__shift_9__pad_1);

  $dumpvars(0,shifter_right_tc__width_6__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_6__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_6__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_6__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_6__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_6__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_6__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_6__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_6__shift_8__pad_0);

  $dumpvars(0,shifter_right_tc__width_6__shift_9__pad_0);

  $dumpvars(0,shifter_right_tc__width_6__shift_10__pad_0);

  $dumpvars(0,shifter_right_tc__width_6__shift_11__pad_0);

  $dumpvars(0,shifter_right_tc__width_6__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_6__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_6__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_6__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_6__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_6__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_6__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_6__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_6__shift_8__pad_1);

  $dumpvars(0,shifter_right_tc__width_6__shift_9__pad_1);

  $dumpvars(0,shifter_right_tc__width_6__shift_10__pad_1);

  $dumpvars(0,shifter_right_tc__width_6__shift_11__pad_1);

  $dumpvars(0,shifter_right_tc__width_7__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_7__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_7__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_7__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_7__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_7__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_7__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_7__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_7__shift_8__pad_0);

  $dumpvars(0,shifter_right_tc__width_7__shift_9__pad_0);

  $dumpvars(0,shifter_right_tc__width_7__shift_10__pad_0);

  $dumpvars(0,shifter_right_tc__width_7__shift_11__pad_0);

  $dumpvars(0,shifter_right_tc__width_7__shift_12__pad_0);

  $dumpvars(0,shifter_right_tc__width_7__shift_13__pad_0);

  $dumpvars(0,shifter_right_tc__width_7__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_7__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_7__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_7__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_7__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_7__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_7__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_7__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_7__shift_8__pad_1);

  $dumpvars(0,shifter_right_tc__width_7__shift_9__pad_1);

  $dumpvars(0,shifter_right_tc__width_7__shift_10__pad_1);

  $dumpvars(0,shifter_right_tc__width_7__shift_11__pad_1);

  $dumpvars(0,shifter_right_tc__width_7__shift_12__pad_1);

  $dumpvars(0,shifter_right_tc__width_7__shift_13__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_8__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_9__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_10__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_11__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_12__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_13__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_14__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_15__pad_0);

  $dumpvars(0,shifter_right_tc__width_8__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_8__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_9__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_10__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_11__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_12__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_13__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_14__pad_1);

  $dumpvars(0,shifter_right_tc__width_8__shift_15__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_8__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_9__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_10__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_11__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_12__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_13__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_14__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_15__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_16__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_17__pad_0);

  $dumpvars(0,shifter_right_tc__width_9__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_8__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_9__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_10__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_11__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_12__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_13__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_14__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_15__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_16__pad_1);

  $dumpvars(0,shifter_right_tc__width_9__shift_17__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_8__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_9__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_10__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_11__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_12__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_13__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_14__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_15__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_16__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_17__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_18__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_19__pad_0);

  $dumpvars(0,shifter_right_tc__width_10__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_8__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_9__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_10__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_11__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_12__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_13__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_14__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_15__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_16__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_17__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_18__pad_1);

  $dumpvars(0,shifter_right_tc__width_10__shift_19__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_8__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_9__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_10__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_11__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_12__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_13__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_14__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_15__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_16__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_17__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_18__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_19__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_20__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_21__pad_0);

  $dumpvars(0,shifter_right_tc__width_11__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_8__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_9__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_10__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_11__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_12__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_13__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_14__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_15__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_16__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_17__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_18__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_19__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_20__pad_1);

  $dumpvars(0,shifter_right_tc__width_11__shift_21__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_8__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_9__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_10__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_11__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_12__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_13__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_14__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_15__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_16__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_17__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_18__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_19__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_20__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_21__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_22__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_23__pad_0);

  $dumpvars(0,shifter_right_tc__width_12__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_8__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_9__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_10__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_11__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_12__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_13__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_14__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_15__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_16__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_17__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_18__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_19__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_20__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_21__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_22__pad_1);

  $dumpvars(0,shifter_right_tc__width_12__shift_23__pad_1);

  $dumpvars(0,shifter_right_tc__width_16__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_16__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_16__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_16__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_16__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_16__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_16__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_16__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_16__shift_8__pad_0);

  $dumpvars(0,shifter_right_tc__width_16__shift_15__pad_0);

  $dumpvars(0,shifter_right_tc__width_16__shift_16__pad_0);

  $dumpvars(0,shifter_right_tc__width_16__shift_17__pad_0);

  $dumpvars(0,shifter_right_tc__width_16__shift_24__pad_0);

  $dumpvars(0,shifter_right_tc__width_16__shift_31__pad_0);

  $dumpvars(0,shifter_right_tc__width_16__shift_32__pad_0);

  $dumpvars(0,shifter_right_tc__width_16__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_16__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_16__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_16__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_16__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_16__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_16__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_16__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_16__shift_8__pad_1);

  $dumpvars(0,shifter_right_tc__width_16__shift_15__pad_1);

  $dumpvars(0,shifter_right_tc__width_16__shift_16__pad_1);

  $dumpvars(0,shifter_right_tc__width_16__shift_17__pad_1);

  $dumpvars(0,shifter_right_tc__width_16__shift_24__pad_1);

  $dumpvars(0,shifter_right_tc__width_16__shift_31__pad_1);

  $dumpvars(0,shifter_right_tc__width_16__shift_32__pad_1);

  $dumpvars(0,shifter_right_tc__width_24__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_24__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_24__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_24__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_24__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_24__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_24__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_24__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_24__shift_12__pad_0);

  $dumpvars(0,shifter_right_tc__width_24__shift_23__pad_0);

  $dumpvars(0,shifter_right_tc__width_24__shift_24__pad_0);

  $dumpvars(0,shifter_right_tc__width_24__shift_25__pad_0);

  $dumpvars(0,shifter_right_tc__width_24__shift_36__pad_0);

  $dumpvars(0,shifter_right_tc__width_24__shift_47__pad_0);

  $dumpvars(0,shifter_right_tc__width_24__shift_48__pad_0);

  $dumpvars(0,shifter_right_tc__width_24__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_24__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_24__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_24__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_24__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_24__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_24__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_24__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_24__shift_12__pad_1);

  $dumpvars(0,shifter_right_tc__width_24__shift_23__pad_1);

  $dumpvars(0,shifter_right_tc__width_24__shift_24__pad_1);

  $dumpvars(0,shifter_right_tc__width_24__shift_25__pad_1);

  $dumpvars(0,shifter_right_tc__width_24__shift_36__pad_1);

  $dumpvars(0,shifter_right_tc__width_24__shift_47__pad_1);

  $dumpvars(0,shifter_right_tc__width_24__shift_48__pad_1);

  $dumpvars(0,shifter_right_tc__width_32__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_32__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_32__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_32__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_32__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_32__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_32__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_32__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_32__shift_16__pad_0);

  $dumpvars(0,shifter_right_tc__width_32__shift_31__pad_0);

  $dumpvars(0,shifter_right_tc__width_32__shift_32__pad_0);

  $dumpvars(0,shifter_right_tc__width_32__shift_33__pad_0);

  $dumpvars(0,shifter_right_tc__width_32__shift_48__pad_0);

  $dumpvars(0,shifter_right_tc__width_32__shift_63__pad_0);

  $dumpvars(0,shifter_right_tc__width_32__shift_64__pad_0);

  $dumpvars(0,shifter_right_tc__width_32__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_32__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_32__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_32__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_32__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_32__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_32__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_32__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_32__shift_16__pad_1);

  $dumpvars(0,shifter_right_tc__width_32__shift_31__pad_1);

  $dumpvars(0,shifter_right_tc__width_32__shift_32__pad_1);

  $dumpvars(0,shifter_right_tc__width_32__shift_33__pad_1);

  $dumpvars(0,shifter_right_tc__width_32__shift_48__pad_1);

  $dumpvars(0,shifter_right_tc__width_32__shift_63__pad_1);

  $dumpvars(0,shifter_right_tc__width_32__shift_64__pad_1);

  $dumpvars(0,shifter_right_tc__width_48__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_48__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_48__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_48__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_48__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_48__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_48__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_48__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_48__shift_24__pad_0);

  $dumpvars(0,shifter_right_tc__width_48__shift_47__pad_0);

  $dumpvars(0,shifter_right_tc__width_48__shift_48__pad_0);

  $dumpvars(0,shifter_right_tc__width_48__shift_49__pad_0);

  $dumpvars(0,shifter_right_tc__width_48__shift_72__pad_0);

  $dumpvars(0,shifter_right_tc__width_48__shift_95__pad_0);

  $dumpvars(0,shifter_right_tc__width_48__shift_96__pad_0);

  $dumpvars(0,shifter_right_tc__width_48__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_48__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_48__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_48__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_48__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_48__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_48__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_48__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_48__shift_24__pad_1);

  $dumpvars(0,shifter_right_tc__width_48__shift_47__pad_1);

  $dumpvars(0,shifter_right_tc__width_48__shift_48__pad_1);

  $dumpvars(0,shifter_right_tc__width_48__shift_49__pad_1);

  $dumpvars(0,shifter_right_tc__width_48__shift_72__pad_1);

  $dumpvars(0,shifter_right_tc__width_48__shift_95__pad_1);

  $dumpvars(0,shifter_right_tc__width_48__shift_96__pad_1);

  $dumpvars(0,shifter_right_tc__width_64__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_64__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_64__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_64__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_64__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_64__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_64__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_64__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_64__shift_32__pad_0);

  $dumpvars(0,shifter_right_tc__width_64__shift_63__pad_0);

  $dumpvars(0,shifter_right_tc__width_64__shift_64__pad_0);

  $dumpvars(0,shifter_right_tc__width_64__shift_65__pad_0);

  $dumpvars(0,shifter_right_tc__width_64__shift_96__pad_0);

  $dumpvars(0,shifter_right_tc__width_64__shift_127__pad_0);

  $dumpvars(0,shifter_right_tc__width_64__shift_128__pad_0);

  $dumpvars(0,shifter_right_tc__width_64__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_64__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_64__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_64__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_64__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_64__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_64__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_64__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_64__shift_32__pad_1);

  $dumpvars(0,shifter_right_tc__width_64__shift_63__pad_1);

  $dumpvars(0,shifter_right_tc__width_64__shift_64__pad_1);

  $dumpvars(0,shifter_right_tc__width_64__shift_65__pad_1);

  $dumpvars(0,shifter_right_tc__width_64__shift_96__pad_1);

  $dumpvars(0,shifter_right_tc__width_64__shift_127__pad_1);

  $dumpvars(0,shifter_right_tc__width_64__shift_128__pad_1);

  $dumpvars(0,shifter_right_tc__width_128__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_128__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_128__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_128__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_128__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_128__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_128__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_128__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_128__shift_64__pad_0);

  $dumpvars(0,shifter_right_tc__width_128__shift_127__pad_0);

  $dumpvars(0,shifter_right_tc__width_128__shift_128__pad_0);

  $dumpvars(0,shifter_right_tc__width_128__shift_129__pad_0);

  $dumpvars(0,shifter_right_tc__width_128__shift_192__pad_0);

  $dumpvars(0,shifter_right_tc__width_128__shift_255__pad_0);

  $dumpvars(0,shifter_right_tc__width_128__shift_256__pad_0);

  $dumpvars(0,shifter_right_tc__width_128__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_128__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_128__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_128__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_128__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_128__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_128__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_128__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_128__shift_64__pad_1);

  $dumpvars(0,shifter_right_tc__width_128__shift_127__pad_1);

  $dumpvars(0,shifter_right_tc__width_128__shift_128__pad_1);

  $dumpvars(0,shifter_right_tc__width_128__shift_129__pad_1);

  $dumpvars(0,shifter_right_tc__width_128__shift_192__pad_1);

  $dumpvars(0,shifter_right_tc__width_128__shift_255__pad_1);

  $dumpvars(0,shifter_right_tc__width_128__shift_256__pad_1);

  $dumpvars(0,shifter_right_tc__width_256__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_256__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_256__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_256__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_256__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_256__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_256__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_256__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_256__shift_128__pad_0);

  $dumpvars(0,shifter_right_tc__width_256__shift_255__pad_0);

  $dumpvars(0,shifter_right_tc__width_256__shift_256__pad_0);

  $dumpvars(0,shifter_right_tc__width_256__shift_257__pad_0);

  $dumpvars(0,shifter_right_tc__width_256__shift_384__pad_0);

  $dumpvars(0,shifter_right_tc__width_256__shift_511__pad_0);

  $dumpvars(0,shifter_right_tc__width_256__shift_512__pad_0);

  $dumpvars(0,shifter_right_tc__width_256__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_256__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_256__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_256__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_256__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_256__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_256__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_256__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_256__shift_128__pad_1);

  $dumpvars(0,shifter_right_tc__width_256__shift_255__pad_1);

  $dumpvars(0,shifter_right_tc__width_256__shift_256__pad_1);

  $dumpvars(0,shifter_right_tc__width_256__shift_257__pad_1);

  $dumpvars(0,shifter_right_tc__width_256__shift_384__pad_1);

  $dumpvars(0,shifter_right_tc__width_256__shift_511__pad_1);

  $dumpvars(0,shifter_right_tc__width_256__shift_512__pad_1);

  $dumpvars(0,shifter_right_tc__width_512__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_512__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_512__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_512__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_512__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_512__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_512__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_512__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_512__shift_256__pad_0);

  $dumpvars(0,shifter_right_tc__width_512__shift_511__pad_0);

  $dumpvars(0,shifter_right_tc__width_512__shift_512__pad_0);

  $dumpvars(0,shifter_right_tc__width_512__shift_513__pad_0);

  $dumpvars(0,shifter_right_tc__width_512__shift_768__pad_0);

  $dumpvars(0,shifter_right_tc__width_512__shift_1023__pad_0);

  $dumpvars(0,shifter_right_tc__width_512__shift_1024__pad_0);

  $dumpvars(0,shifter_right_tc__width_512__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_512__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_512__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_512__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_512__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_512__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_512__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_512__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_512__shift_256__pad_1);

  $dumpvars(0,shifter_right_tc__width_512__shift_511__pad_1);

  $dumpvars(0,shifter_right_tc__width_512__shift_512__pad_1);

  $dumpvars(0,shifter_right_tc__width_512__shift_513__pad_1);

  $dumpvars(0,shifter_right_tc__width_512__shift_768__pad_1);

  $dumpvars(0,shifter_right_tc__width_512__shift_1023__pad_1);

  $dumpvars(0,shifter_right_tc__width_512__shift_1024__pad_1);

  $dumpvars(0,shifter_right_tc__width_1024__shift_0__pad_0);

  $dumpvars(0,shifter_right_tc__width_1024__shift_1__pad_0);

  $dumpvars(0,shifter_right_tc__width_1024__shift_2__pad_0);

  $dumpvars(0,shifter_right_tc__width_1024__shift_3__pad_0);

  $dumpvars(0,shifter_right_tc__width_1024__shift_4__pad_0);

  $dumpvars(0,shifter_right_tc__width_1024__shift_5__pad_0);

  $dumpvars(0,shifter_right_tc__width_1024__shift_6__pad_0);

  $dumpvars(0,shifter_right_tc__width_1024__shift_7__pad_0);

  $dumpvars(0,shifter_right_tc__width_1024__shift_512__pad_0);

  $dumpvars(0,shifter_right_tc__width_1024__shift_1023__pad_0);

  $dumpvars(0,shifter_right_tc__width_1024__shift_1024__pad_0);

  $dumpvars(0,shifter_right_tc__width_1024__shift_1025__pad_0);

  $dumpvars(0,shifter_right_tc__width_1024__shift_1536__pad_0);

  $dumpvars(0,shifter_right_tc__width_1024__shift_2047__pad_0);

  $dumpvars(0,shifter_right_tc__width_1024__shift_2048__pad_0);

  $dumpvars(0,shifter_right_tc__width_1024__shift_0__pad_1);

  $dumpvars(0,shifter_right_tc__width_1024__shift_1__pad_1);

  $dumpvars(0,shifter_right_tc__width_1024__shift_2__pad_1);

  $dumpvars(0,shifter_right_tc__width_1024__shift_3__pad_1);

  $dumpvars(0,shifter_right_tc__width_1024__shift_4__pad_1);

  $dumpvars(0,shifter_right_tc__width_1024__shift_5__pad_1);

  $dumpvars(0,shifter_right_tc__width_1024__shift_6__pad_1);

  $dumpvars(0,shifter_right_tc__width_1024__shift_7__pad_1);

  $dumpvars(0,shifter_right_tc__width_1024__shift_512__pad_1);

  $dumpvars(0,shifter_right_tc__width_1024__shift_1023__pad_1);

  $dumpvars(0,shifter_right_tc__width_1024__shift_1024__pad_1);

  $dumpvars(0,shifter_right_tc__width_1024__shift_1025__pad_1);

  $dumpvars(0,shifter_right_tc__width_1024__shift_1536__pad_1);

  $dumpvars(0,shifter_right_tc__width_1024__shift_2047__pad_1);

  $dumpvars(0,shifter_right_tc__width_1024__shift_2048__pad_1);


  // Initialization


  start__shifter_right_tc__width_1__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_1__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_1__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_1__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_2__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_2__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_2__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_2__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_2__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_2__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_2__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_2__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_3__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_3__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_3__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_3__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_3__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_3__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_3__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_3__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_3__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_3__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_3__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_3__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_4__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_4__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_4__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_4__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_4__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_4__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_4__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_4__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_4__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_4__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_4__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_4__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_4__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_4__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_4__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_4__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_5__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_5__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_5__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_5__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_5__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_5__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_5__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_5__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_5__shift_8__pad_0 = 0;

  start__shifter_right_tc__width_5__shift_9__pad_0 = 0;

  start__shifter_right_tc__width_5__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_5__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_5__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_5__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_5__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_5__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_5__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_5__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_5__shift_8__pad_1 = 0;

  start__shifter_right_tc__width_5__shift_9__pad_1 = 0;

  start__shifter_right_tc__width_6__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_6__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_6__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_6__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_6__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_6__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_6__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_6__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_6__shift_8__pad_0 = 0;

  start__shifter_right_tc__width_6__shift_9__pad_0 = 0;

  start__shifter_right_tc__width_6__shift_10__pad_0 = 0;

  start__shifter_right_tc__width_6__shift_11__pad_0 = 0;

  start__shifter_right_tc__width_6__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_6__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_6__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_6__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_6__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_6__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_6__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_6__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_6__shift_8__pad_1 = 0;

  start__shifter_right_tc__width_6__shift_9__pad_1 = 0;

  start__shifter_right_tc__width_6__shift_10__pad_1 = 0;

  start__shifter_right_tc__width_6__shift_11__pad_1 = 0;

  start__shifter_right_tc__width_7__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_7__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_7__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_7__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_7__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_7__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_7__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_7__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_7__shift_8__pad_0 = 0;

  start__shifter_right_tc__width_7__shift_9__pad_0 = 0;

  start__shifter_right_tc__width_7__shift_10__pad_0 = 0;

  start__shifter_right_tc__width_7__shift_11__pad_0 = 0;

  start__shifter_right_tc__width_7__shift_12__pad_0 = 0;

  start__shifter_right_tc__width_7__shift_13__pad_0 = 0;

  start__shifter_right_tc__width_7__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_7__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_7__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_7__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_7__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_7__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_7__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_7__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_7__shift_8__pad_1 = 0;

  start__shifter_right_tc__width_7__shift_9__pad_1 = 0;

  start__shifter_right_tc__width_7__shift_10__pad_1 = 0;

  start__shifter_right_tc__width_7__shift_11__pad_1 = 0;

  start__shifter_right_tc__width_7__shift_12__pad_1 = 0;

  start__shifter_right_tc__width_7__shift_13__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_8__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_9__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_10__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_11__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_12__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_13__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_14__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_15__pad_0 = 0;

  start__shifter_right_tc__width_8__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_8__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_9__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_10__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_11__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_12__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_13__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_14__pad_1 = 0;

  start__shifter_right_tc__width_8__shift_15__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_8__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_9__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_10__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_11__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_12__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_13__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_14__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_15__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_16__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_17__pad_0 = 0;

  start__shifter_right_tc__width_9__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_8__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_9__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_10__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_11__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_12__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_13__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_14__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_15__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_16__pad_1 = 0;

  start__shifter_right_tc__width_9__shift_17__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_8__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_9__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_10__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_11__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_12__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_13__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_14__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_15__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_16__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_17__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_18__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_19__pad_0 = 0;

  start__shifter_right_tc__width_10__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_8__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_9__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_10__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_11__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_12__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_13__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_14__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_15__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_16__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_17__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_18__pad_1 = 0;

  start__shifter_right_tc__width_10__shift_19__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_8__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_9__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_10__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_11__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_12__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_13__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_14__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_15__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_16__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_17__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_18__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_19__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_20__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_21__pad_0 = 0;

  start__shifter_right_tc__width_11__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_8__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_9__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_10__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_11__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_12__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_13__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_14__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_15__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_16__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_17__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_18__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_19__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_20__pad_1 = 0;

  start__shifter_right_tc__width_11__shift_21__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_8__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_9__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_10__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_11__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_12__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_13__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_14__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_15__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_16__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_17__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_18__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_19__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_20__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_21__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_22__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_23__pad_0 = 0;

  start__shifter_right_tc__width_12__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_8__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_9__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_10__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_11__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_12__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_13__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_14__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_15__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_16__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_17__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_18__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_19__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_20__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_21__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_22__pad_1 = 0;

  start__shifter_right_tc__width_12__shift_23__pad_1 = 0;

  start__shifter_right_tc__width_16__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_16__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_16__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_16__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_16__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_16__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_16__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_16__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_16__shift_8__pad_0 = 0;

  start__shifter_right_tc__width_16__shift_15__pad_0 = 0;

  start__shifter_right_tc__width_16__shift_16__pad_0 = 0;

  start__shifter_right_tc__width_16__shift_17__pad_0 = 0;

  start__shifter_right_tc__width_16__shift_24__pad_0 = 0;

  start__shifter_right_tc__width_16__shift_31__pad_0 = 0;

  start__shifter_right_tc__width_16__shift_32__pad_0 = 0;

  start__shifter_right_tc__width_16__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_16__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_16__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_16__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_16__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_16__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_16__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_16__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_16__shift_8__pad_1 = 0;

  start__shifter_right_tc__width_16__shift_15__pad_1 = 0;

  start__shifter_right_tc__width_16__shift_16__pad_1 = 0;

  start__shifter_right_tc__width_16__shift_17__pad_1 = 0;

  start__shifter_right_tc__width_16__shift_24__pad_1 = 0;

  start__shifter_right_tc__width_16__shift_31__pad_1 = 0;

  start__shifter_right_tc__width_16__shift_32__pad_1 = 0;

  start__shifter_right_tc__width_24__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_24__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_24__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_24__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_24__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_24__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_24__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_24__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_24__shift_12__pad_0 = 0;

  start__shifter_right_tc__width_24__shift_23__pad_0 = 0;

  start__shifter_right_tc__width_24__shift_24__pad_0 = 0;

  start__shifter_right_tc__width_24__shift_25__pad_0 = 0;

  start__shifter_right_tc__width_24__shift_36__pad_0 = 0;

  start__shifter_right_tc__width_24__shift_47__pad_0 = 0;

  start__shifter_right_tc__width_24__shift_48__pad_0 = 0;

  start__shifter_right_tc__width_24__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_24__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_24__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_24__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_24__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_24__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_24__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_24__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_24__shift_12__pad_1 = 0;

  start__shifter_right_tc__width_24__shift_23__pad_1 = 0;

  start__shifter_right_tc__width_24__shift_24__pad_1 = 0;

  start__shifter_right_tc__width_24__shift_25__pad_1 = 0;

  start__shifter_right_tc__width_24__shift_36__pad_1 = 0;

  start__shifter_right_tc__width_24__shift_47__pad_1 = 0;

  start__shifter_right_tc__width_24__shift_48__pad_1 = 0;

  start__shifter_right_tc__width_32__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_32__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_32__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_32__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_32__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_32__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_32__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_32__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_32__shift_16__pad_0 = 0;

  start__shifter_right_tc__width_32__shift_31__pad_0 = 0;

  start__shifter_right_tc__width_32__shift_32__pad_0 = 0;

  start__shifter_right_tc__width_32__shift_33__pad_0 = 0;

  start__shifter_right_tc__width_32__shift_48__pad_0 = 0;

  start__shifter_right_tc__width_32__shift_63__pad_0 = 0;

  start__shifter_right_tc__width_32__shift_64__pad_0 = 0;

  start__shifter_right_tc__width_32__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_32__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_32__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_32__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_32__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_32__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_32__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_32__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_32__shift_16__pad_1 = 0;

  start__shifter_right_tc__width_32__shift_31__pad_1 = 0;

  start__shifter_right_tc__width_32__shift_32__pad_1 = 0;

  start__shifter_right_tc__width_32__shift_33__pad_1 = 0;

  start__shifter_right_tc__width_32__shift_48__pad_1 = 0;

  start__shifter_right_tc__width_32__shift_63__pad_1 = 0;

  start__shifter_right_tc__width_32__shift_64__pad_1 = 0;

  start__shifter_right_tc__width_48__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_48__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_48__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_48__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_48__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_48__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_48__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_48__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_48__shift_24__pad_0 = 0;

  start__shifter_right_tc__width_48__shift_47__pad_0 = 0;

  start__shifter_right_tc__width_48__shift_48__pad_0 = 0;

  start__shifter_right_tc__width_48__shift_49__pad_0 = 0;

  start__shifter_right_tc__width_48__shift_72__pad_0 = 0;

  start__shifter_right_tc__width_48__shift_95__pad_0 = 0;

  start__shifter_right_tc__width_48__shift_96__pad_0 = 0;

  start__shifter_right_tc__width_48__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_48__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_48__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_48__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_48__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_48__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_48__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_48__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_48__shift_24__pad_1 = 0;

  start__shifter_right_tc__width_48__shift_47__pad_1 = 0;

  start__shifter_right_tc__width_48__shift_48__pad_1 = 0;

  start__shifter_right_tc__width_48__shift_49__pad_1 = 0;

  start__shifter_right_tc__width_48__shift_72__pad_1 = 0;

  start__shifter_right_tc__width_48__shift_95__pad_1 = 0;

  start__shifter_right_tc__width_48__shift_96__pad_1 = 0;

  start__shifter_right_tc__width_64__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_64__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_64__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_64__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_64__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_64__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_64__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_64__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_64__shift_32__pad_0 = 0;

  start__shifter_right_tc__width_64__shift_63__pad_0 = 0;

  start__shifter_right_tc__width_64__shift_64__pad_0 = 0;

  start__shifter_right_tc__width_64__shift_65__pad_0 = 0;

  start__shifter_right_tc__width_64__shift_96__pad_0 = 0;

  start__shifter_right_tc__width_64__shift_127__pad_0 = 0;

  start__shifter_right_tc__width_64__shift_128__pad_0 = 0;

  start__shifter_right_tc__width_64__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_64__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_64__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_64__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_64__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_64__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_64__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_64__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_64__shift_32__pad_1 = 0;

  start__shifter_right_tc__width_64__shift_63__pad_1 = 0;

  start__shifter_right_tc__width_64__shift_64__pad_1 = 0;

  start__shifter_right_tc__width_64__shift_65__pad_1 = 0;

  start__shifter_right_tc__width_64__shift_96__pad_1 = 0;

  start__shifter_right_tc__width_64__shift_127__pad_1 = 0;

  start__shifter_right_tc__width_64__shift_128__pad_1 = 0;

  start__shifter_right_tc__width_128__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_128__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_128__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_128__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_128__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_128__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_128__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_128__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_128__shift_64__pad_0 = 0;

  start__shifter_right_tc__width_128__shift_127__pad_0 = 0;

  start__shifter_right_tc__width_128__shift_128__pad_0 = 0;

  start__shifter_right_tc__width_128__shift_129__pad_0 = 0;

  start__shifter_right_tc__width_128__shift_192__pad_0 = 0;

  start__shifter_right_tc__width_128__shift_255__pad_0 = 0;

  start__shifter_right_tc__width_128__shift_256__pad_0 = 0;

  start__shifter_right_tc__width_128__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_128__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_128__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_128__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_128__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_128__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_128__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_128__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_128__shift_64__pad_1 = 0;

  start__shifter_right_tc__width_128__shift_127__pad_1 = 0;

  start__shifter_right_tc__width_128__shift_128__pad_1 = 0;

  start__shifter_right_tc__width_128__shift_129__pad_1 = 0;

  start__shifter_right_tc__width_128__shift_192__pad_1 = 0;

  start__shifter_right_tc__width_128__shift_255__pad_1 = 0;

  start__shifter_right_tc__width_128__shift_256__pad_1 = 0;

  start__shifter_right_tc__width_256__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_256__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_256__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_256__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_256__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_256__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_256__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_256__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_256__shift_128__pad_0 = 0;

  start__shifter_right_tc__width_256__shift_255__pad_0 = 0;

  start__shifter_right_tc__width_256__shift_256__pad_0 = 0;

  start__shifter_right_tc__width_256__shift_257__pad_0 = 0;

  start__shifter_right_tc__width_256__shift_384__pad_0 = 0;

  start__shifter_right_tc__width_256__shift_511__pad_0 = 0;

  start__shifter_right_tc__width_256__shift_512__pad_0 = 0;

  start__shifter_right_tc__width_256__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_256__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_256__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_256__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_256__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_256__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_256__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_256__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_256__shift_128__pad_1 = 0;

  start__shifter_right_tc__width_256__shift_255__pad_1 = 0;

  start__shifter_right_tc__width_256__shift_256__pad_1 = 0;

  start__shifter_right_tc__width_256__shift_257__pad_1 = 0;

  start__shifter_right_tc__width_256__shift_384__pad_1 = 0;

  start__shifter_right_tc__width_256__shift_511__pad_1 = 0;

  start__shifter_right_tc__width_256__shift_512__pad_1 = 0;

  start__shifter_right_tc__width_512__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_512__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_512__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_512__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_512__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_512__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_512__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_512__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_512__shift_256__pad_0 = 0;

  start__shifter_right_tc__width_512__shift_511__pad_0 = 0;

  start__shifter_right_tc__width_512__shift_512__pad_0 = 0;

  start__shifter_right_tc__width_512__shift_513__pad_0 = 0;

  start__shifter_right_tc__width_512__shift_768__pad_0 = 0;

  start__shifter_right_tc__width_512__shift_1023__pad_0 = 0;

  start__shifter_right_tc__width_512__shift_1024__pad_0 = 0;

  start__shifter_right_tc__width_512__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_512__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_512__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_512__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_512__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_512__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_512__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_512__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_512__shift_256__pad_1 = 0;

  start__shifter_right_tc__width_512__shift_511__pad_1 = 0;

  start__shifter_right_tc__width_512__shift_512__pad_1 = 0;

  start__shifter_right_tc__width_512__shift_513__pad_1 = 0;

  start__shifter_right_tc__width_512__shift_768__pad_1 = 0;

  start__shifter_right_tc__width_512__shift_1023__pad_1 = 0;

  start__shifter_right_tc__width_512__shift_1024__pad_1 = 0;

  start__shifter_right_tc__width_1024__shift_0__pad_0 = 0;

  start__shifter_right_tc__width_1024__shift_1__pad_0 = 0;

  start__shifter_right_tc__width_1024__shift_2__pad_0 = 0;

  start__shifter_right_tc__width_1024__shift_3__pad_0 = 0;

  start__shifter_right_tc__width_1024__shift_4__pad_0 = 0;

  start__shifter_right_tc__width_1024__shift_5__pad_0 = 0;

  start__shifter_right_tc__width_1024__shift_6__pad_0 = 0;

  start__shifter_right_tc__width_1024__shift_7__pad_0 = 0;

  start__shifter_right_tc__width_1024__shift_512__pad_0 = 0;

  start__shifter_right_tc__width_1024__shift_1023__pad_0 = 0;

  start__shifter_right_tc__width_1024__shift_1024__pad_0 = 0;

  start__shifter_right_tc__width_1024__shift_1025__pad_0 = 0;

  start__shifter_right_tc__width_1024__shift_1536__pad_0 = 0;

  start__shifter_right_tc__width_1024__shift_2047__pad_0 = 0;

  start__shifter_right_tc__width_1024__shift_2048__pad_0 = 0;

  start__shifter_right_tc__width_1024__shift_0__pad_1 = 0;

  start__shifter_right_tc__width_1024__shift_1__pad_1 = 0;

  start__shifter_right_tc__width_1024__shift_2__pad_1 = 0;

  start__shifter_right_tc__width_1024__shift_3__pad_1 = 0;

  start__shifter_right_tc__width_1024__shift_4__pad_1 = 0;

  start__shifter_right_tc__width_1024__shift_5__pad_1 = 0;

  start__shifter_right_tc__width_1024__shift_6__pad_1 = 0;

  start__shifter_right_tc__width_1024__shift_7__pad_1 = 0;

  start__shifter_right_tc__width_1024__shift_512__pad_1 = 0;

  start__shifter_right_tc__width_1024__shift_1023__pad_1 = 0;

  start__shifter_right_tc__width_1024__shift_1024__pad_1 = 0;

  start__shifter_right_tc__width_1024__shift_1025__pad_1 = 0;

  start__shifter_right_tc__width_1024__shift_1536__pad_1 = 0;

  start__shifter_right_tc__width_1024__shift_2047__pad_1 = 0;

  start__shifter_right_tc__width_1024__shift_2048__pad_1 = 0;


  // Start testbenches

  start__shifter_right_tc__width_1__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_1__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_1__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_1__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_1__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_1__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_1__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_1__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_2__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_2__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_2__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_2__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_2__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_2__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_2__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_2__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_2__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_2__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_2__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_2__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_2__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_2__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_2__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_2__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_3__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_3__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_3__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_3__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_3__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_3__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_3__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_3__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_3__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_3__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_3__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_3__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_3__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_3__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_3__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_3__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_3__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_3__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_3__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_3__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_3__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_3__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_3__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_3__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_4__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_4__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_4__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_4__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_4__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_4__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_4__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_4__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_4__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_4__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_4__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_4__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_4__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_4__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_4__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_4__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_4__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_4__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_4__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_4__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_4__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_4__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_4__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_4__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_4__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_4__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_4__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_4__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_4__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_4__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_4__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_4__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_5__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_5__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_5__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_5__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_5__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_5__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_5__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_5__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_5__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_5__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_5__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_5__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_5__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_5__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_5__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_5__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_5__shift_8__pad_0 = 1;
  while(!shifter_right_tc__width_5__shift_8__pad_0.finished) #(1);

  start__shifter_right_tc__width_5__shift_9__pad_0 = 1;
  while(!shifter_right_tc__width_5__shift_9__pad_0.finished) #(1);

  start__shifter_right_tc__width_5__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_5__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_5__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_5__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_5__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_5__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_5__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_5__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_5__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_5__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_5__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_5__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_5__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_5__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_5__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_5__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_5__shift_8__pad_1 = 1;
  while(!shifter_right_tc__width_5__shift_8__pad_1.finished) #(1);

  start__shifter_right_tc__width_5__shift_9__pad_1 = 1;
  while(!shifter_right_tc__width_5__shift_9__pad_1.finished) #(1);

  start__shifter_right_tc__width_6__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_6__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_6__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_6__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_6__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_6__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_6__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_6__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_6__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_6__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_6__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_6__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_6__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_6__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_6__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_6__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_6__shift_8__pad_0 = 1;
  while(!shifter_right_tc__width_6__shift_8__pad_0.finished) #(1);

  start__shifter_right_tc__width_6__shift_9__pad_0 = 1;
  while(!shifter_right_tc__width_6__shift_9__pad_0.finished) #(1);

  start__shifter_right_tc__width_6__shift_10__pad_0 = 1;
  while(!shifter_right_tc__width_6__shift_10__pad_0.finished) #(1);

  start__shifter_right_tc__width_6__shift_11__pad_0 = 1;
  while(!shifter_right_tc__width_6__shift_11__pad_0.finished) #(1);

  start__shifter_right_tc__width_6__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_6__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_6__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_6__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_6__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_6__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_6__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_6__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_6__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_6__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_6__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_6__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_6__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_6__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_6__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_6__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_6__shift_8__pad_1 = 1;
  while(!shifter_right_tc__width_6__shift_8__pad_1.finished) #(1);

  start__shifter_right_tc__width_6__shift_9__pad_1 = 1;
  while(!shifter_right_tc__width_6__shift_9__pad_1.finished) #(1);

  start__shifter_right_tc__width_6__shift_10__pad_1 = 1;
  while(!shifter_right_tc__width_6__shift_10__pad_1.finished) #(1);

  start__shifter_right_tc__width_6__shift_11__pad_1 = 1;
  while(!shifter_right_tc__width_6__shift_11__pad_1.finished) #(1);

  start__shifter_right_tc__width_7__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_7__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_7__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_7__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_7__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_7__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_7__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_7__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_7__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_7__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_7__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_7__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_7__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_7__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_7__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_7__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_7__shift_8__pad_0 = 1;
  while(!shifter_right_tc__width_7__shift_8__pad_0.finished) #(1);

  start__shifter_right_tc__width_7__shift_9__pad_0 = 1;
  while(!shifter_right_tc__width_7__shift_9__pad_0.finished) #(1);

  start__shifter_right_tc__width_7__shift_10__pad_0 = 1;
  while(!shifter_right_tc__width_7__shift_10__pad_0.finished) #(1);

  start__shifter_right_tc__width_7__shift_11__pad_0 = 1;
  while(!shifter_right_tc__width_7__shift_11__pad_0.finished) #(1);

  start__shifter_right_tc__width_7__shift_12__pad_0 = 1;
  while(!shifter_right_tc__width_7__shift_12__pad_0.finished) #(1);

  start__shifter_right_tc__width_7__shift_13__pad_0 = 1;
  while(!shifter_right_tc__width_7__shift_13__pad_0.finished) #(1);

  start__shifter_right_tc__width_7__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_7__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_7__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_7__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_7__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_7__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_7__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_7__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_7__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_7__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_7__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_7__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_7__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_7__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_7__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_7__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_7__shift_8__pad_1 = 1;
  while(!shifter_right_tc__width_7__shift_8__pad_1.finished) #(1);

  start__shifter_right_tc__width_7__shift_9__pad_1 = 1;
  while(!shifter_right_tc__width_7__shift_9__pad_1.finished) #(1);

  start__shifter_right_tc__width_7__shift_10__pad_1 = 1;
  while(!shifter_right_tc__width_7__shift_10__pad_1.finished) #(1);

  start__shifter_right_tc__width_7__shift_11__pad_1 = 1;
  while(!shifter_right_tc__width_7__shift_11__pad_1.finished) #(1);

  start__shifter_right_tc__width_7__shift_12__pad_1 = 1;
  while(!shifter_right_tc__width_7__shift_12__pad_1.finished) #(1);

  start__shifter_right_tc__width_7__shift_13__pad_1 = 1;
  while(!shifter_right_tc__width_7__shift_13__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_8__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_8__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_9__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_9__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_10__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_10__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_11__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_11__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_12__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_12__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_13__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_13__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_14__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_14__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_15__pad_0 = 1;
  while(!shifter_right_tc__width_8__shift_15__pad_0.finished) #(1);

  start__shifter_right_tc__width_8__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_8__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_8__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_9__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_9__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_10__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_10__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_11__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_11__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_12__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_12__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_13__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_13__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_14__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_14__pad_1.finished) #(1);

  start__shifter_right_tc__width_8__shift_15__pad_1 = 1;
  while(!shifter_right_tc__width_8__shift_15__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_8__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_8__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_9__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_9__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_10__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_10__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_11__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_11__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_12__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_12__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_13__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_13__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_14__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_14__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_15__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_15__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_16__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_16__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_17__pad_0 = 1;
  while(!shifter_right_tc__width_9__shift_17__pad_0.finished) #(1);

  start__shifter_right_tc__width_9__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_8__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_8__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_9__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_9__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_10__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_10__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_11__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_11__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_12__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_12__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_13__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_13__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_14__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_14__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_15__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_15__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_16__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_16__pad_1.finished) #(1);

  start__shifter_right_tc__width_9__shift_17__pad_1 = 1;
  while(!shifter_right_tc__width_9__shift_17__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_8__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_8__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_9__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_9__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_10__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_10__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_11__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_11__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_12__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_12__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_13__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_13__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_14__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_14__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_15__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_15__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_16__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_16__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_17__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_17__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_18__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_18__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_19__pad_0 = 1;
  while(!shifter_right_tc__width_10__shift_19__pad_0.finished) #(1);

  start__shifter_right_tc__width_10__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_8__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_8__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_9__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_9__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_10__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_10__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_11__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_11__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_12__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_12__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_13__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_13__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_14__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_14__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_15__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_15__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_16__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_16__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_17__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_17__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_18__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_18__pad_1.finished) #(1);

  start__shifter_right_tc__width_10__shift_19__pad_1 = 1;
  while(!shifter_right_tc__width_10__shift_19__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_8__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_8__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_9__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_9__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_10__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_10__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_11__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_11__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_12__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_12__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_13__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_13__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_14__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_14__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_15__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_15__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_16__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_16__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_17__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_17__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_18__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_18__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_19__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_19__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_20__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_20__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_21__pad_0 = 1;
  while(!shifter_right_tc__width_11__shift_21__pad_0.finished) #(1);

  start__shifter_right_tc__width_11__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_8__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_8__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_9__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_9__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_10__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_10__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_11__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_11__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_12__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_12__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_13__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_13__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_14__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_14__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_15__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_15__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_16__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_16__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_17__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_17__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_18__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_18__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_19__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_19__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_20__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_20__pad_1.finished) #(1);

  start__shifter_right_tc__width_11__shift_21__pad_1 = 1;
  while(!shifter_right_tc__width_11__shift_21__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_8__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_8__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_9__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_9__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_10__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_10__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_11__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_11__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_12__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_12__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_13__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_13__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_14__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_14__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_15__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_15__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_16__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_16__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_17__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_17__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_18__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_18__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_19__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_19__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_20__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_20__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_21__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_21__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_22__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_22__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_23__pad_0 = 1;
  while(!shifter_right_tc__width_12__shift_23__pad_0.finished) #(1);

  start__shifter_right_tc__width_12__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_8__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_8__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_9__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_9__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_10__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_10__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_11__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_11__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_12__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_12__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_13__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_13__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_14__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_14__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_15__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_15__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_16__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_16__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_17__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_17__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_18__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_18__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_19__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_19__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_20__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_20__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_21__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_21__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_22__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_22__pad_1.finished) #(1);

  start__shifter_right_tc__width_12__shift_23__pad_1 = 1;
  while(!shifter_right_tc__width_12__shift_23__pad_1.finished) #(1);

  start__shifter_right_tc__width_16__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_16__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_16__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_16__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_16__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_16__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_16__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_16__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_16__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_16__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_16__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_16__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_16__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_16__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_16__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_16__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_16__shift_8__pad_0 = 1;
  while(!shifter_right_tc__width_16__shift_8__pad_0.finished) #(1);

  start__shifter_right_tc__width_16__shift_15__pad_0 = 1;
  while(!shifter_right_tc__width_16__shift_15__pad_0.finished) #(1);

  start__shifter_right_tc__width_16__shift_16__pad_0 = 1;
  while(!shifter_right_tc__width_16__shift_16__pad_0.finished) #(1);

  start__shifter_right_tc__width_16__shift_17__pad_0 = 1;
  while(!shifter_right_tc__width_16__shift_17__pad_0.finished) #(1);

  start__shifter_right_tc__width_16__shift_24__pad_0 = 1;
  while(!shifter_right_tc__width_16__shift_24__pad_0.finished) #(1);

  start__shifter_right_tc__width_16__shift_31__pad_0 = 1;
  while(!shifter_right_tc__width_16__shift_31__pad_0.finished) #(1);

  start__shifter_right_tc__width_16__shift_32__pad_0 = 1;
  while(!shifter_right_tc__width_16__shift_32__pad_0.finished) #(1);

  start__shifter_right_tc__width_16__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_16__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_16__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_16__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_16__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_16__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_16__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_16__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_16__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_16__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_16__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_16__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_16__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_16__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_16__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_16__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_16__shift_8__pad_1 = 1;
  while(!shifter_right_tc__width_16__shift_8__pad_1.finished) #(1);

  start__shifter_right_tc__width_16__shift_15__pad_1 = 1;
  while(!shifter_right_tc__width_16__shift_15__pad_1.finished) #(1);

  start__shifter_right_tc__width_16__shift_16__pad_1 = 1;
  while(!shifter_right_tc__width_16__shift_16__pad_1.finished) #(1);

  start__shifter_right_tc__width_16__shift_17__pad_1 = 1;
  while(!shifter_right_tc__width_16__shift_17__pad_1.finished) #(1);

  start__shifter_right_tc__width_16__shift_24__pad_1 = 1;
  while(!shifter_right_tc__width_16__shift_24__pad_1.finished) #(1);

  start__shifter_right_tc__width_16__shift_31__pad_1 = 1;
  while(!shifter_right_tc__width_16__shift_31__pad_1.finished) #(1);

  start__shifter_right_tc__width_16__shift_32__pad_1 = 1;
  while(!shifter_right_tc__width_16__shift_32__pad_1.finished) #(1);

  start__shifter_right_tc__width_24__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_24__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_24__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_24__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_24__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_24__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_24__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_24__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_24__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_24__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_24__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_24__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_24__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_24__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_24__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_24__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_24__shift_12__pad_0 = 1;
  while(!shifter_right_tc__width_24__shift_12__pad_0.finished) #(1);

  start__shifter_right_tc__width_24__shift_23__pad_0 = 1;
  while(!shifter_right_tc__width_24__shift_23__pad_0.finished) #(1);

  start__shifter_right_tc__width_24__shift_24__pad_0 = 1;
  while(!shifter_right_tc__width_24__shift_24__pad_0.finished) #(1);

  start__shifter_right_tc__width_24__shift_25__pad_0 = 1;
  while(!shifter_right_tc__width_24__shift_25__pad_0.finished) #(1);

  start__shifter_right_tc__width_24__shift_36__pad_0 = 1;
  while(!shifter_right_tc__width_24__shift_36__pad_0.finished) #(1);

  start__shifter_right_tc__width_24__shift_47__pad_0 = 1;
  while(!shifter_right_tc__width_24__shift_47__pad_0.finished) #(1);

  start__shifter_right_tc__width_24__shift_48__pad_0 = 1;
  while(!shifter_right_tc__width_24__shift_48__pad_0.finished) #(1);

  start__shifter_right_tc__width_24__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_24__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_24__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_24__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_24__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_24__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_24__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_24__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_24__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_24__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_24__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_24__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_24__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_24__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_24__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_24__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_24__shift_12__pad_1 = 1;
  while(!shifter_right_tc__width_24__shift_12__pad_1.finished) #(1);

  start__shifter_right_tc__width_24__shift_23__pad_1 = 1;
  while(!shifter_right_tc__width_24__shift_23__pad_1.finished) #(1);

  start__shifter_right_tc__width_24__shift_24__pad_1 = 1;
  while(!shifter_right_tc__width_24__shift_24__pad_1.finished) #(1);

  start__shifter_right_tc__width_24__shift_25__pad_1 = 1;
  while(!shifter_right_tc__width_24__shift_25__pad_1.finished) #(1);

  start__shifter_right_tc__width_24__shift_36__pad_1 = 1;
  while(!shifter_right_tc__width_24__shift_36__pad_1.finished) #(1);

  start__shifter_right_tc__width_24__shift_47__pad_1 = 1;
  while(!shifter_right_tc__width_24__shift_47__pad_1.finished) #(1);

  start__shifter_right_tc__width_24__shift_48__pad_1 = 1;
  while(!shifter_right_tc__width_24__shift_48__pad_1.finished) #(1);

  start__shifter_right_tc__width_32__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_32__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_32__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_32__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_32__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_32__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_32__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_32__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_32__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_32__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_32__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_32__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_32__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_32__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_32__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_32__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_32__shift_16__pad_0 = 1;
  while(!shifter_right_tc__width_32__shift_16__pad_0.finished) #(1);

  start__shifter_right_tc__width_32__shift_31__pad_0 = 1;
  while(!shifter_right_tc__width_32__shift_31__pad_0.finished) #(1);

  start__shifter_right_tc__width_32__shift_32__pad_0 = 1;
  while(!shifter_right_tc__width_32__shift_32__pad_0.finished) #(1);

  start__shifter_right_tc__width_32__shift_33__pad_0 = 1;
  while(!shifter_right_tc__width_32__shift_33__pad_0.finished) #(1);

  start__shifter_right_tc__width_32__shift_48__pad_0 = 1;
  while(!shifter_right_tc__width_32__shift_48__pad_0.finished) #(1);

  start__shifter_right_tc__width_32__shift_63__pad_0 = 1;
  while(!shifter_right_tc__width_32__shift_63__pad_0.finished) #(1);

  start__shifter_right_tc__width_32__shift_64__pad_0 = 1;
  while(!shifter_right_tc__width_32__shift_64__pad_0.finished) #(1);

  start__shifter_right_tc__width_32__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_32__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_32__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_32__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_32__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_32__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_32__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_32__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_32__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_32__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_32__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_32__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_32__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_32__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_32__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_32__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_32__shift_16__pad_1 = 1;
  while(!shifter_right_tc__width_32__shift_16__pad_1.finished) #(1);

  start__shifter_right_tc__width_32__shift_31__pad_1 = 1;
  while(!shifter_right_tc__width_32__shift_31__pad_1.finished) #(1);

  start__shifter_right_tc__width_32__shift_32__pad_1 = 1;
  while(!shifter_right_tc__width_32__shift_32__pad_1.finished) #(1);

  start__shifter_right_tc__width_32__shift_33__pad_1 = 1;
  while(!shifter_right_tc__width_32__shift_33__pad_1.finished) #(1);

  start__shifter_right_tc__width_32__shift_48__pad_1 = 1;
  while(!shifter_right_tc__width_32__shift_48__pad_1.finished) #(1);

  start__shifter_right_tc__width_32__shift_63__pad_1 = 1;
  while(!shifter_right_tc__width_32__shift_63__pad_1.finished) #(1);

  start__shifter_right_tc__width_32__shift_64__pad_1 = 1;
  while(!shifter_right_tc__width_32__shift_64__pad_1.finished) #(1);

  start__shifter_right_tc__width_48__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_48__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_48__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_48__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_48__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_48__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_48__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_48__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_48__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_48__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_48__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_48__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_48__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_48__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_48__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_48__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_48__shift_24__pad_0 = 1;
  while(!shifter_right_tc__width_48__shift_24__pad_0.finished) #(1);

  start__shifter_right_tc__width_48__shift_47__pad_0 = 1;
  while(!shifter_right_tc__width_48__shift_47__pad_0.finished) #(1);

  start__shifter_right_tc__width_48__shift_48__pad_0 = 1;
  while(!shifter_right_tc__width_48__shift_48__pad_0.finished) #(1);

  start__shifter_right_tc__width_48__shift_49__pad_0 = 1;
  while(!shifter_right_tc__width_48__shift_49__pad_0.finished) #(1);

  start__shifter_right_tc__width_48__shift_72__pad_0 = 1;
  while(!shifter_right_tc__width_48__shift_72__pad_0.finished) #(1);

  start__shifter_right_tc__width_48__shift_95__pad_0 = 1;
  while(!shifter_right_tc__width_48__shift_95__pad_0.finished) #(1);

  start__shifter_right_tc__width_48__shift_96__pad_0 = 1;
  while(!shifter_right_tc__width_48__shift_96__pad_0.finished) #(1);

  start__shifter_right_tc__width_48__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_48__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_48__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_48__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_48__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_48__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_48__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_48__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_48__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_48__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_48__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_48__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_48__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_48__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_48__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_48__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_48__shift_24__pad_1 = 1;
  while(!shifter_right_tc__width_48__shift_24__pad_1.finished) #(1);

  start__shifter_right_tc__width_48__shift_47__pad_1 = 1;
  while(!shifter_right_tc__width_48__shift_47__pad_1.finished) #(1);

  start__shifter_right_tc__width_48__shift_48__pad_1 = 1;
  while(!shifter_right_tc__width_48__shift_48__pad_1.finished) #(1);

  start__shifter_right_tc__width_48__shift_49__pad_1 = 1;
  while(!shifter_right_tc__width_48__shift_49__pad_1.finished) #(1);

  start__shifter_right_tc__width_48__shift_72__pad_1 = 1;
  while(!shifter_right_tc__width_48__shift_72__pad_1.finished) #(1);

  start__shifter_right_tc__width_48__shift_95__pad_1 = 1;
  while(!shifter_right_tc__width_48__shift_95__pad_1.finished) #(1);

  start__shifter_right_tc__width_48__shift_96__pad_1 = 1;
  while(!shifter_right_tc__width_48__shift_96__pad_1.finished) #(1);

  start__shifter_right_tc__width_64__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_64__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_64__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_64__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_64__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_64__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_64__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_64__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_64__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_64__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_64__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_64__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_64__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_64__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_64__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_64__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_64__shift_32__pad_0 = 1;
  while(!shifter_right_tc__width_64__shift_32__pad_0.finished) #(1);

  start__shifter_right_tc__width_64__shift_63__pad_0 = 1;
  while(!shifter_right_tc__width_64__shift_63__pad_0.finished) #(1);

  start__shifter_right_tc__width_64__shift_64__pad_0 = 1;
  while(!shifter_right_tc__width_64__shift_64__pad_0.finished) #(1);

  start__shifter_right_tc__width_64__shift_65__pad_0 = 1;
  while(!shifter_right_tc__width_64__shift_65__pad_0.finished) #(1);

  start__shifter_right_tc__width_64__shift_96__pad_0 = 1;
  while(!shifter_right_tc__width_64__shift_96__pad_0.finished) #(1);

  start__shifter_right_tc__width_64__shift_127__pad_0 = 1;
  while(!shifter_right_tc__width_64__shift_127__pad_0.finished) #(1);

  start__shifter_right_tc__width_64__shift_128__pad_0 = 1;
  while(!shifter_right_tc__width_64__shift_128__pad_0.finished) #(1);

  start__shifter_right_tc__width_64__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_64__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_64__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_64__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_64__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_64__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_64__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_64__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_64__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_64__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_64__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_64__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_64__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_64__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_64__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_64__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_64__shift_32__pad_1 = 1;
  while(!shifter_right_tc__width_64__shift_32__pad_1.finished) #(1);

  start__shifter_right_tc__width_64__shift_63__pad_1 = 1;
  while(!shifter_right_tc__width_64__shift_63__pad_1.finished) #(1);

  start__shifter_right_tc__width_64__shift_64__pad_1 = 1;
  while(!shifter_right_tc__width_64__shift_64__pad_1.finished) #(1);

  start__shifter_right_tc__width_64__shift_65__pad_1 = 1;
  while(!shifter_right_tc__width_64__shift_65__pad_1.finished) #(1);

  start__shifter_right_tc__width_64__shift_96__pad_1 = 1;
  while(!shifter_right_tc__width_64__shift_96__pad_1.finished) #(1);

  start__shifter_right_tc__width_64__shift_127__pad_1 = 1;
  while(!shifter_right_tc__width_64__shift_127__pad_1.finished) #(1);

  start__shifter_right_tc__width_64__shift_128__pad_1 = 1;
  while(!shifter_right_tc__width_64__shift_128__pad_1.finished) #(1);

  start__shifter_right_tc__width_128__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_128__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_128__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_128__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_128__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_128__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_128__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_128__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_128__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_128__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_128__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_128__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_128__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_128__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_128__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_128__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_128__shift_64__pad_0 = 1;
  while(!shifter_right_tc__width_128__shift_64__pad_0.finished) #(1);

  start__shifter_right_tc__width_128__shift_127__pad_0 = 1;
  while(!shifter_right_tc__width_128__shift_127__pad_0.finished) #(1);

  start__shifter_right_tc__width_128__shift_128__pad_0 = 1;
  while(!shifter_right_tc__width_128__shift_128__pad_0.finished) #(1);

  start__shifter_right_tc__width_128__shift_129__pad_0 = 1;
  while(!shifter_right_tc__width_128__shift_129__pad_0.finished) #(1);

  start__shifter_right_tc__width_128__shift_192__pad_0 = 1;
  while(!shifter_right_tc__width_128__shift_192__pad_0.finished) #(1);

  start__shifter_right_tc__width_128__shift_255__pad_0 = 1;
  while(!shifter_right_tc__width_128__shift_255__pad_0.finished) #(1);

  start__shifter_right_tc__width_128__shift_256__pad_0 = 1;
  while(!shifter_right_tc__width_128__shift_256__pad_0.finished) #(1);

  start__shifter_right_tc__width_128__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_128__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_128__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_128__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_128__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_128__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_128__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_128__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_128__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_128__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_128__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_128__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_128__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_128__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_128__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_128__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_128__shift_64__pad_1 = 1;
  while(!shifter_right_tc__width_128__shift_64__pad_1.finished) #(1);

  start__shifter_right_tc__width_128__shift_127__pad_1 = 1;
  while(!shifter_right_tc__width_128__shift_127__pad_1.finished) #(1);

  start__shifter_right_tc__width_128__shift_128__pad_1 = 1;
  while(!shifter_right_tc__width_128__shift_128__pad_1.finished) #(1);

  start__shifter_right_tc__width_128__shift_129__pad_1 = 1;
  while(!shifter_right_tc__width_128__shift_129__pad_1.finished) #(1);

  start__shifter_right_tc__width_128__shift_192__pad_1 = 1;
  while(!shifter_right_tc__width_128__shift_192__pad_1.finished) #(1);

  start__shifter_right_tc__width_128__shift_255__pad_1 = 1;
  while(!shifter_right_tc__width_128__shift_255__pad_1.finished) #(1);

  start__shifter_right_tc__width_128__shift_256__pad_1 = 1;
  while(!shifter_right_tc__width_128__shift_256__pad_1.finished) #(1);

  start__shifter_right_tc__width_256__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_256__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_256__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_256__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_256__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_256__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_256__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_256__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_256__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_256__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_256__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_256__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_256__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_256__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_256__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_256__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_256__shift_128__pad_0 = 1;
  while(!shifter_right_tc__width_256__shift_128__pad_0.finished) #(1);

  start__shifter_right_tc__width_256__shift_255__pad_0 = 1;
  while(!shifter_right_tc__width_256__shift_255__pad_0.finished) #(1);

  start__shifter_right_tc__width_256__shift_256__pad_0 = 1;
  while(!shifter_right_tc__width_256__shift_256__pad_0.finished) #(1);

  start__shifter_right_tc__width_256__shift_257__pad_0 = 1;
  while(!shifter_right_tc__width_256__shift_257__pad_0.finished) #(1);

  start__shifter_right_tc__width_256__shift_384__pad_0 = 1;
  while(!shifter_right_tc__width_256__shift_384__pad_0.finished) #(1);

  start__shifter_right_tc__width_256__shift_511__pad_0 = 1;
  while(!shifter_right_tc__width_256__shift_511__pad_0.finished) #(1);

  start__shifter_right_tc__width_256__shift_512__pad_0 = 1;
  while(!shifter_right_tc__width_256__shift_512__pad_0.finished) #(1);

  start__shifter_right_tc__width_256__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_256__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_256__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_256__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_256__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_256__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_256__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_256__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_256__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_256__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_256__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_256__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_256__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_256__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_256__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_256__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_256__shift_128__pad_1 = 1;
  while(!shifter_right_tc__width_256__shift_128__pad_1.finished) #(1);

  start__shifter_right_tc__width_256__shift_255__pad_1 = 1;
  while(!shifter_right_tc__width_256__shift_255__pad_1.finished) #(1);

  start__shifter_right_tc__width_256__shift_256__pad_1 = 1;
  while(!shifter_right_tc__width_256__shift_256__pad_1.finished) #(1);

  start__shifter_right_tc__width_256__shift_257__pad_1 = 1;
  while(!shifter_right_tc__width_256__shift_257__pad_1.finished) #(1);

  start__shifter_right_tc__width_256__shift_384__pad_1 = 1;
  while(!shifter_right_tc__width_256__shift_384__pad_1.finished) #(1);

  start__shifter_right_tc__width_256__shift_511__pad_1 = 1;
  while(!shifter_right_tc__width_256__shift_511__pad_1.finished) #(1);

  start__shifter_right_tc__width_256__shift_512__pad_1 = 1;
  while(!shifter_right_tc__width_256__shift_512__pad_1.finished) #(1);

  start__shifter_right_tc__width_512__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_512__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_512__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_512__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_512__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_512__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_512__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_512__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_512__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_512__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_512__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_512__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_512__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_512__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_512__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_512__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_512__shift_256__pad_0 = 1;
  while(!shifter_right_tc__width_512__shift_256__pad_0.finished) #(1);

  start__shifter_right_tc__width_512__shift_511__pad_0 = 1;
  while(!shifter_right_tc__width_512__shift_511__pad_0.finished) #(1);

  start__shifter_right_tc__width_512__shift_512__pad_0 = 1;
  while(!shifter_right_tc__width_512__shift_512__pad_0.finished) #(1);

  start__shifter_right_tc__width_512__shift_513__pad_0 = 1;
  while(!shifter_right_tc__width_512__shift_513__pad_0.finished) #(1);

  start__shifter_right_tc__width_512__shift_768__pad_0 = 1;
  while(!shifter_right_tc__width_512__shift_768__pad_0.finished) #(1);

  start__shifter_right_tc__width_512__shift_1023__pad_0 = 1;
  while(!shifter_right_tc__width_512__shift_1023__pad_0.finished) #(1);

  start__shifter_right_tc__width_512__shift_1024__pad_0 = 1;
  while(!shifter_right_tc__width_512__shift_1024__pad_0.finished) #(1);

  start__shifter_right_tc__width_512__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_512__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_512__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_512__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_512__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_512__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_512__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_512__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_512__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_512__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_512__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_512__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_512__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_512__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_512__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_512__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_512__shift_256__pad_1 = 1;
  while(!shifter_right_tc__width_512__shift_256__pad_1.finished) #(1);

  start__shifter_right_tc__width_512__shift_511__pad_1 = 1;
  while(!shifter_right_tc__width_512__shift_511__pad_1.finished) #(1);

  start__shifter_right_tc__width_512__shift_512__pad_1 = 1;
  while(!shifter_right_tc__width_512__shift_512__pad_1.finished) #(1);

  start__shifter_right_tc__width_512__shift_513__pad_1 = 1;
  while(!shifter_right_tc__width_512__shift_513__pad_1.finished) #(1);

  start__shifter_right_tc__width_512__shift_768__pad_1 = 1;
  while(!shifter_right_tc__width_512__shift_768__pad_1.finished) #(1);

  start__shifter_right_tc__width_512__shift_1023__pad_1 = 1;
  while(!shifter_right_tc__width_512__shift_1023__pad_1.finished) #(1);

  start__shifter_right_tc__width_512__shift_1024__pad_1 = 1;
  while(!shifter_right_tc__width_512__shift_1024__pad_1.finished) #(1);

  start__shifter_right_tc__width_1024__shift_0__pad_0 = 1;
  while(!shifter_right_tc__width_1024__shift_0__pad_0.finished) #(1);

  start__shifter_right_tc__width_1024__shift_1__pad_0 = 1;
  while(!shifter_right_tc__width_1024__shift_1__pad_0.finished) #(1);

  start__shifter_right_tc__width_1024__shift_2__pad_0 = 1;
  while(!shifter_right_tc__width_1024__shift_2__pad_0.finished) #(1);

  start__shifter_right_tc__width_1024__shift_3__pad_0 = 1;
  while(!shifter_right_tc__width_1024__shift_3__pad_0.finished) #(1);

  start__shifter_right_tc__width_1024__shift_4__pad_0 = 1;
  while(!shifter_right_tc__width_1024__shift_4__pad_0.finished) #(1);

  start__shifter_right_tc__width_1024__shift_5__pad_0 = 1;
  while(!shifter_right_tc__width_1024__shift_5__pad_0.finished) #(1);

  start__shifter_right_tc__width_1024__shift_6__pad_0 = 1;
  while(!shifter_right_tc__width_1024__shift_6__pad_0.finished) #(1);

  start__shifter_right_tc__width_1024__shift_7__pad_0 = 1;
  while(!shifter_right_tc__width_1024__shift_7__pad_0.finished) #(1);

  start__shifter_right_tc__width_1024__shift_512__pad_0 = 1;
  while(!shifter_right_tc__width_1024__shift_512__pad_0.finished) #(1);

  start__shifter_right_tc__width_1024__shift_1023__pad_0 = 1;
  while(!shifter_right_tc__width_1024__shift_1023__pad_0.finished) #(1);

  start__shifter_right_tc__width_1024__shift_1024__pad_0 = 1;
  while(!shifter_right_tc__width_1024__shift_1024__pad_0.finished) #(1);

  start__shifter_right_tc__width_1024__shift_1025__pad_0 = 1;
  while(!shifter_right_tc__width_1024__shift_1025__pad_0.finished) #(1);

  start__shifter_right_tc__width_1024__shift_1536__pad_0 = 1;
  while(!shifter_right_tc__width_1024__shift_1536__pad_0.finished) #(1);

  start__shifter_right_tc__width_1024__shift_2047__pad_0 = 1;
  while(!shifter_right_tc__width_1024__shift_2047__pad_0.finished) #(1);

  start__shifter_right_tc__width_1024__shift_2048__pad_0 = 1;
  while(!shifter_right_tc__width_1024__shift_2048__pad_0.finished) #(1);

  start__shifter_right_tc__width_1024__shift_0__pad_1 = 1;
  while(!shifter_right_tc__width_1024__shift_0__pad_1.finished) #(1);

  start__shifter_right_tc__width_1024__shift_1__pad_1 = 1;
  while(!shifter_right_tc__width_1024__shift_1__pad_1.finished) #(1);

  start__shifter_right_tc__width_1024__shift_2__pad_1 = 1;
  while(!shifter_right_tc__width_1024__shift_2__pad_1.finished) #(1);

  start__shifter_right_tc__width_1024__shift_3__pad_1 = 1;
  while(!shifter_right_tc__width_1024__shift_3__pad_1.finished) #(1);

  start__shifter_right_tc__width_1024__shift_4__pad_1 = 1;
  while(!shifter_right_tc__width_1024__shift_4__pad_1.finished) #(1);

  start__shifter_right_tc__width_1024__shift_5__pad_1 = 1;
  while(!shifter_right_tc__width_1024__shift_5__pad_1.finished) #(1);

  start__shifter_right_tc__width_1024__shift_6__pad_1 = 1;
  while(!shifter_right_tc__width_1024__shift_6__pad_1.finished) #(1);

  start__shifter_right_tc__width_1024__shift_7__pad_1 = 1;
  while(!shifter_right_tc__width_1024__shift_7__pad_1.finished) #(1);

  start__shifter_right_tc__width_1024__shift_512__pad_1 = 1;
  while(!shifter_right_tc__width_1024__shift_512__pad_1.finished) #(1);

  start__shifter_right_tc__width_1024__shift_1023__pad_1 = 1;
  while(!shifter_right_tc__width_1024__shift_1023__pad_1.finished) #(1);

  start__shifter_right_tc__width_1024__shift_1024__pad_1 = 1;
  while(!shifter_right_tc__width_1024__shift_1024__pad_1.finished) #(1);

  start__shifter_right_tc__width_1024__shift_1025__pad_1 = 1;
  while(!shifter_right_tc__width_1024__shift_1025__pad_1.finished) #(1);

  start__shifter_right_tc__width_1024__shift_1536__pad_1 = 1;
  while(!shifter_right_tc__width_1024__shift_1536__pad_1.finished) #(1);

  start__shifter_right_tc__width_1024__shift_2047__pad_1 = 1;
  while(!shifter_right_tc__width_1024__shift_2047__pad_1.finished) #(1);

  start__shifter_right_tc__width_1024__shift_2048__pad_1 = 1;
  while(!shifter_right_tc__width_1024__shift_2048__pad_1.finished) #(1);


  // Finish
  $finish();
end

endmodule