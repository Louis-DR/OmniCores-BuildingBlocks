`include "hamming.svh"

`ifndef GET_EXTENDED_HAMMING_PARITY_WIDTH
`define GET_EXTENDED_HAMMING_PARITY_WIDTH(DATA_WIDTH) \
  (DATA_WIDTH <= 65519) ? `GET_HAMMING_PARITY_WIDTH(DATA_WIDTH) + 1 : -1
`endif

`ifndef GET_EXTENDED_HAMMING_DATA_WIDTH
`define GET_EXTENDED_HAMMING_DATA_WIDTH(PARITY_WIDTH) \
  (PARITY_WIDTH <= 17) ? `GET_HAMMING_DATA_WIDTH(PARITY_WIDTH-1) : -1
`endif

`ifndef GET_EXTENDED_HAMMING_PARITY_WIDTH_FROM_BLOCK_WIDTH
`define GET_EXTENDED_HAMMING_PARITY_WIDTH_FROM_BLOCK_WIDTH(BLOCK_WIDTH) \
  (BLOCK_WIDTH <= 65536) ? `GET_HAMMING_PARITY_WIDTH_FROM_BLOCK_WIDTH(BLOCK_WIDTH-1) + 1 : -1
`endif

`ifndef GET_EXTENDED_HAMMING_DATA_WIDTH_FROM_BLOCK_WIDTH
`define GET_EXTENDED_HAMMING_DATA_WIDTH_FROM_BLOCK_WIDTH(BLOCK_WIDTH) \
  (BLOCK_WIDTH <= 65536) ? `GET_HAMMING_DATA_WIDTH_FROM_BLOCK_WIDTH(BLOCK_WIDTH-1) - 1 : -1
`endif

`ifndef GET_EXTENDED_HAMMING_UPPER_BLOCK_WIDTH
`define GET_EXTENDED_HAMMING_UPPER_BLOCK_WIDTH(BLOCK_WIDTH) \
  (BLOCK_WIDTH <= 65536) ? `GET_HAMMING_UPPER_BLOCK_WIDTH(BLOCK_WIDTH-1) + 1 : -1
`endif
