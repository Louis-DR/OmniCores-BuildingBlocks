
`ifndef INFINITE
`define INFINITE (1/0)
`endif

typedef bit bool;

localparam bool true  = 1'b1;
localparam bool false = 1'b0;
