// ╔═══════════════════════════════════════════════════════════════════════════╗
// ║ Project:     OmniCores-BuildingBlocks                                     ║
// ║ Author:      Louis Duret-Robert - louisduret@gmail.com                    ║
// ║ Website:     louis-dr.github.io                                           ║
// ║ License:     MIT License                                                  ║
// ║ File:        extended_hamming_checker.sv                                  ║
// ╟───────────────────────────────────────────────────────────────────────────╢
// ║ Description: Detects correctable single-bit errors and uncorrectable      ║
// ║              double-bit errors in data with extended Hamming code.        ║
// ║                                                                           ║
// ╚═══════════════════════════════════════════════════════════════════════════╝



`include "extended_hamming.svh"



module extended_hamming_checker #(
  parameter  DATA_WIDTH   = 8,
  localparam PARITY_WIDTH = `GET_EXTENDED_HAMMING_PARITY_WIDTH(DATA_WIDTH),
  localparam BLOCK_WIDTH  = DATA_WIDTH + PARITY_WIDTH
) (
  input   [DATA_WIDTH-1:0] data,
  input [PARITY_WIDTH-1:0] code,
  output                   correctable_error,
  output                   uncorrectable_error
);

// Pad the data to the message length corresponding to the number of parity bits
localparam PADDED_DATA_WIDTH = `GET_EXTENDED_HAMMING_DATA_WIDTH(PARITY_WIDTH);
logic [PADDED_DATA_WIDTH-1:0] data_padded;
assign data_padded = {{(PADDED_DATA_WIDTH - DATA_WIDTH){1'b0}}, data};

// Pad the block
localparam PADDED_BLOCK_WIDTH = PADDED_DATA_WIDTH + PARITY_WIDTH;
logic [PADDED_BLOCK_WIDTH-1:0] block_padded;

extended_hamming_block_packer #(
  .DATA_WIDTH ( PADDED_DATA_WIDTH )
) packager (
  .data  ( data_padded  ),
  .code  ( code         ),
  .block ( block_padded )
);

extended_hamming_block_checker #(
  .BLOCK_WIDTH ( PADDED_BLOCK_WIDTH )
) block_checker (
  .block               ( block_padded        ),
  .correctable_error   ( correctable_error   ),
  .uncorrectable_error ( uncorrectable_error )
);

endmodule