// ╔═══════════════════════════════════════════════════════════════════════════╗
// ║ Project:     OmniCores-BuildingBlocks                                     ║
// ║ Author:      Louis Duret-Robert - louisduret@gmail.com                    ║
// ║ Website:     louis-dr.github.io                                           ║
// ║ License:     MIT License                                                  ║
// ║ File:        rotator_left.tb.sv                                           ║
// ╟───────────────────────────────────────────────────────────────────────────╢
// ║ This file is generated from the template rotator_left.tb.sv.j2 by J2GPP.  ║
// ║ Do not edit it directly.                                                  ║
// ╟───────────────────────────────────────────────────────────────────────────╢
// ║ Description: Top-level testbench for the static left rotator.             ║
// ║                                                                           ║
// ╚═══════════════════════════════════════════════════════════════════════════╝



`timescale 1ns/1ns



module rotator_left_tb ();


logic start__rotator_left_tc__width_1__rotation_0;
logic start__rotator_left_tc__width_1__rotation_1;

logic start__rotator_left_tc__width_2__rotation_0;
logic start__rotator_left_tc__width_2__rotation_1;
logic start__rotator_left_tc__width_2__rotation_2;
logic start__rotator_left_tc__width_2__rotation_3;

logic start__rotator_left_tc__width_3__rotation_0;
logic start__rotator_left_tc__width_3__rotation_1;
logic start__rotator_left_tc__width_3__rotation_2;
logic start__rotator_left_tc__width_3__rotation_3;
logic start__rotator_left_tc__width_3__rotation_4;
logic start__rotator_left_tc__width_3__rotation_5;

logic start__rotator_left_tc__width_4__rotation_0;
logic start__rotator_left_tc__width_4__rotation_1;
logic start__rotator_left_tc__width_4__rotation_2;
logic start__rotator_left_tc__width_4__rotation_3;
logic start__rotator_left_tc__width_4__rotation_4;
logic start__rotator_left_tc__width_4__rotation_5;
logic start__rotator_left_tc__width_4__rotation_6;
logic start__rotator_left_tc__width_4__rotation_7;

logic start__rotator_left_tc__width_5__rotation_0;
logic start__rotator_left_tc__width_5__rotation_1;
logic start__rotator_left_tc__width_5__rotation_2;
logic start__rotator_left_tc__width_5__rotation_3;
logic start__rotator_left_tc__width_5__rotation_4;
logic start__rotator_left_tc__width_5__rotation_5;
logic start__rotator_left_tc__width_5__rotation_6;
logic start__rotator_left_tc__width_5__rotation_7;
logic start__rotator_left_tc__width_5__rotation_8;
logic start__rotator_left_tc__width_5__rotation_9;

logic start__rotator_left_tc__width_6__rotation_0;
logic start__rotator_left_tc__width_6__rotation_1;
logic start__rotator_left_tc__width_6__rotation_2;
logic start__rotator_left_tc__width_6__rotation_3;
logic start__rotator_left_tc__width_6__rotation_4;
logic start__rotator_left_tc__width_6__rotation_5;
logic start__rotator_left_tc__width_6__rotation_6;
logic start__rotator_left_tc__width_6__rotation_7;
logic start__rotator_left_tc__width_6__rotation_8;
logic start__rotator_left_tc__width_6__rotation_9;
logic start__rotator_left_tc__width_6__rotation_10;
logic start__rotator_left_tc__width_6__rotation_11;

logic start__rotator_left_tc__width_7__rotation_0;
logic start__rotator_left_tc__width_7__rotation_1;
logic start__rotator_left_tc__width_7__rotation_2;
logic start__rotator_left_tc__width_7__rotation_3;
logic start__rotator_left_tc__width_7__rotation_4;
logic start__rotator_left_tc__width_7__rotation_5;
logic start__rotator_left_tc__width_7__rotation_6;
logic start__rotator_left_tc__width_7__rotation_7;
logic start__rotator_left_tc__width_7__rotation_8;
logic start__rotator_left_tc__width_7__rotation_9;
logic start__rotator_left_tc__width_7__rotation_10;
logic start__rotator_left_tc__width_7__rotation_11;
logic start__rotator_left_tc__width_7__rotation_12;
logic start__rotator_left_tc__width_7__rotation_13;

logic start__rotator_left_tc__width_8__rotation_0;
logic start__rotator_left_tc__width_8__rotation_1;
logic start__rotator_left_tc__width_8__rotation_2;
logic start__rotator_left_tc__width_8__rotation_3;
logic start__rotator_left_tc__width_8__rotation_4;
logic start__rotator_left_tc__width_8__rotation_5;
logic start__rotator_left_tc__width_8__rotation_6;
logic start__rotator_left_tc__width_8__rotation_7;
logic start__rotator_left_tc__width_8__rotation_8;
logic start__rotator_left_tc__width_8__rotation_9;
logic start__rotator_left_tc__width_8__rotation_10;
logic start__rotator_left_tc__width_8__rotation_11;
logic start__rotator_left_tc__width_8__rotation_12;
logic start__rotator_left_tc__width_8__rotation_13;
logic start__rotator_left_tc__width_8__rotation_14;
logic start__rotator_left_tc__width_8__rotation_15;

logic start__rotator_left_tc__width_9__rotation_0;
logic start__rotator_left_tc__width_9__rotation_1;
logic start__rotator_left_tc__width_9__rotation_2;
logic start__rotator_left_tc__width_9__rotation_3;
logic start__rotator_left_tc__width_9__rotation_4;
logic start__rotator_left_tc__width_9__rotation_5;
logic start__rotator_left_tc__width_9__rotation_6;
logic start__rotator_left_tc__width_9__rotation_7;
logic start__rotator_left_tc__width_9__rotation_8;
logic start__rotator_left_tc__width_9__rotation_9;
logic start__rotator_left_tc__width_9__rotation_10;
logic start__rotator_left_tc__width_9__rotation_11;
logic start__rotator_left_tc__width_9__rotation_12;
logic start__rotator_left_tc__width_9__rotation_13;
logic start__rotator_left_tc__width_9__rotation_14;
logic start__rotator_left_tc__width_9__rotation_15;
logic start__rotator_left_tc__width_9__rotation_16;
logic start__rotator_left_tc__width_9__rotation_17;

logic start__rotator_left_tc__width_10__rotation_0;
logic start__rotator_left_tc__width_10__rotation_1;
logic start__rotator_left_tc__width_10__rotation_2;
logic start__rotator_left_tc__width_10__rotation_3;
logic start__rotator_left_tc__width_10__rotation_4;
logic start__rotator_left_tc__width_10__rotation_5;
logic start__rotator_left_tc__width_10__rotation_6;
logic start__rotator_left_tc__width_10__rotation_7;
logic start__rotator_left_tc__width_10__rotation_8;
logic start__rotator_left_tc__width_10__rotation_9;
logic start__rotator_left_tc__width_10__rotation_10;
logic start__rotator_left_tc__width_10__rotation_11;
logic start__rotator_left_tc__width_10__rotation_12;
logic start__rotator_left_tc__width_10__rotation_13;
logic start__rotator_left_tc__width_10__rotation_14;
logic start__rotator_left_tc__width_10__rotation_15;
logic start__rotator_left_tc__width_10__rotation_16;
logic start__rotator_left_tc__width_10__rotation_17;
logic start__rotator_left_tc__width_10__rotation_18;
logic start__rotator_left_tc__width_10__rotation_19;

logic start__rotator_left_tc__width_11__rotation_0;
logic start__rotator_left_tc__width_11__rotation_1;
logic start__rotator_left_tc__width_11__rotation_2;
logic start__rotator_left_tc__width_11__rotation_3;
logic start__rotator_left_tc__width_11__rotation_4;
logic start__rotator_left_tc__width_11__rotation_5;
logic start__rotator_left_tc__width_11__rotation_6;
logic start__rotator_left_tc__width_11__rotation_7;
logic start__rotator_left_tc__width_11__rotation_8;
logic start__rotator_left_tc__width_11__rotation_9;
logic start__rotator_left_tc__width_11__rotation_10;
logic start__rotator_left_tc__width_11__rotation_11;
logic start__rotator_left_tc__width_11__rotation_12;
logic start__rotator_left_tc__width_11__rotation_13;
logic start__rotator_left_tc__width_11__rotation_14;
logic start__rotator_left_tc__width_11__rotation_15;
logic start__rotator_left_tc__width_11__rotation_16;
logic start__rotator_left_tc__width_11__rotation_17;
logic start__rotator_left_tc__width_11__rotation_18;
logic start__rotator_left_tc__width_11__rotation_19;
logic start__rotator_left_tc__width_11__rotation_20;
logic start__rotator_left_tc__width_11__rotation_21;

logic start__rotator_left_tc__width_12__rotation_0;
logic start__rotator_left_tc__width_12__rotation_1;
logic start__rotator_left_tc__width_12__rotation_2;
logic start__rotator_left_tc__width_12__rotation_3;
logic start__rotator_left_tc__width_12__rotation_4;
logic start__rotator_left_tc__width_12__rotation_5;
logic start__rotator_left_tc__width_12__rotation_6;
logic start__rotator_left_tc__width_12__rotation_7;
logic start__rotator_left_tc__width_12__rotation_8;
logic start__rotator_left_tc__width_12__rotation_9;
logic start__rotator_left_tc__width_12__rotation_10;
logic start__rotator_left_tc__width_12__rotation_11;
logic start__rotator_left_tc__width_12__rotation_12;
logic start__rotator_left_tc__width_12__rotation_13;
logic start__rotator_left_tc__width_12__rotation_14;
logic start__rotator_left_tc__width_12__rotation_15;
logic start__rotator_left_tc__width_12__rotation_16;
logic start__rotator_left_tc__width_12__rotation_17;
logic start__rotator_left_tc__width_12__rotation_18;
logic start__rotator_left_tc__width_12__rotation_19;
logic start__rotator_left_tc__width_12__rotation_20;
logic start__rotator_left_tc__width_12__rotation_21;
logic start__rotator_left_tc__width_12__rotation_22;
logic start__rotator_left_tc__width_12__rotation_23;

logic start__rotator_left_tc__width_16__rotation_0;
logic start__rotator_left_tc__width_16__rotation_1;
logic start__rotator_left_tc__width_16__rotation_2;
logic start__rotator_left_tc__width_16__rotation_3;
logic start__rotator_left_tc__width_16__rotation_4;
logic start__rotator_left_tc__width_16__rotation_5;
logic start__rotator_left_tc__width_16__rotation_6;
logic start__rotator_left_tc__width_16__rotation_7;
logic start__rotator_left_tc__width_16__rotation_8;
logic start__rotator_left_tc__width_16__rotation_15;
logic start__rotator_left_tc__width_16__rotation_16;
logic start__rotator_left_tc__width_16__rotation_17;
logic start__rotator_left_tc__width_16__rotation_24;
logic start__rotator_left_tc__width_16__rotation_31;
logic start__rotator_left_tc__width_16__rotation_32;

logic start__rotator_left_tc__width_24__rotation_0;
logic start__rotator_left_tc__width_24__rotation_1;
logic start__rotator_left_tc__width_24__rotation_2;
logic start__rotator_left_tc__width_24__rotation_3;
logic start__rotator_left_tc__width_24__rotation_4;
logic start__rotator_left_tc__width_24__rotation_5;
logic start__rotator_left_tc__width_24__rotation_6;
logic start__rotator_left_tc__width_24__rotation_7;
logic start__rotator_left_tc__width_24__rotation_12;
logic start__rotator_left_tc__width_24__rotation_23;
logic start__rotator_left_tc__width_24__rotation_24;
logic start__rotator_left_tc__width_24__rotation_25;
logic start__rotator_left_tc__width_24__rotation_36;
logic start__rotator_left_tc__width_24__rotation_47;
logic start__rotator_left_tc__width_24__rotation_48;

logic start__rotator_left_tc__width_32__rotation_0;
logic start__rotator_left_tc__width_32__rotation_1;
logic start__rotator_left_tc__width_32__rotation_2;
logic start__rotator_left_tc__width_32__rotation_3;
logic start__rotator_left_tc__width_32__rotation_4;
logic start__rotator_left_tc__width_32__rotation_5;
logic start__rotator_left_tc__width_32__rotation_6;
logic start__rotator_left_tc__width_32__rotation_7;
logic start__rotator_left_tc__width_32__rotation_16;
logic start__rotator_left_tc__width_32__rotation_31;
logic start__rotator_left_tc__width_32__rotation_32;
logic start__rotator_left_tc__width_32__rotation_33;
logic start__rotator_left_tc__width_32__rotation_48;
logic start__rotator_left_tc__width_32__rotation_63;
logic start__rotator_left_tc__width_32__rotation_64;

logic start__rotator_left_tc__width_48__rotation_0;
logic start__rotator_left_tc__width_48__rotation_1;
logic start__rotator_left_tc__width_48__rotation_2;
logic start__rotator_left_tc__width_48__rotation_3;
logic start__rotator_left_tc__width_48__rotation_4;
logic start__rotator_left_tc__width_48__rotation_5;
logic start__rotator_left_tc__width_48__rotation_6;
logic start__rotator_left_tc__width_48__rotation_7;
logic start__rotator_left_tc__width_48__rotation_24;
logic start__rotator_left_tc__width_48__rotation_47;
logic start__rotator_left_tc__width_48__rotation_48;
logic start__rotator_left_tc__width_48__rotation_49;
logic start__rotator_left_tc__width_48__rotation_72;
logic start__rotator_left_tc__width_48__rotation_95;
logic start__rotator_left_tc__width_48__rotation_96;

logic start__rotator_left_tc__width_64__rotation_0;
logic start__rotator_left_tc__width_64__rotation_1;
logic start__rotator_left_tc__width_64__rotation_2;
logic start__rotator_left_tc__width_64__rotation_3;
logic start__rotator_left_tc__width_64__rotation_4;
logic start__rotator_left_tc__width_64__rotation_5;
logic start__rotator_left_tc__width_64__rotation_6;
logic start__rotator_left_tc__width_64__rotation_7;
logic start__rotator_left_tc__width_64__rotation_32;
logic start__rotator_left_tc__width_64__rotation_63;
logic start__rotator_left_tc__width_64__rotation_64;
logic start__rotator_left_tc__width_64__rotation_65;
logic start__rotator_left_tc__width_64__rotation_96;
logic start__rotator_left_tc__width_64__rotation_127;
logic start__rotator_left_tc__width_64__rotation_128;

logic start__rotator_left_tc__width_128__rotation_0;
logic start__rotator_left_tc__width_128__rotation_1;
logic start__rotator_left_tc__width_128__rotation_2;
logic start__rotator_left_tc__width_128__rotation_3;
logic start__rotator_left_tc__width_128__rotation_4;
logic start__rotator_left_tc__width_128__rotation_5;
logic start__rotator_left_tc__width_128__rotation_6;
logic start__rotator_left_tc__width_128__rotation_7;
logic start__rotator_left_tc__width_128__rotation_64;
logic start__rotator_left_tc__width_128__rotation_127;
logic start__rotator_left_tc__width_128__rotation_128;
logic start__rotator_left_tc__width_128__rotation_129;
logic start__rotator_left_tc__width_128__rotation_192;
logic start__rotator_left_tc__width_128__rotation_255;
logic start__rotator_left_tc__width_128__rotation_256;

logic start__rotator_left_tc__width_256__rotation_0;
logic start__rotator_left_tc__width_256__rotation_1;
logic start__rotator_left_tc__width_256__rotation_2;
logic start__rotator_left_tc__width_256__rotation_3;
logic start__rotator_left_tc__width_256__rotation_4;
logic start__rotator_left_tc__width_256__rotation_5;
logic start__rotator_left_tc__width_256__rotation_6;
logic start__rotator_left_tc__width_256__rotation_7;
logic start__rotator_left_tc__width_256__rotation_128;
logic start__rotator_left_tc__width_256__rotation_255;
logic start__rotator_left_tc__width_256__rotation_256;
logic start__rotator_left_tc__width_256__rotation_257;
logic start__rotator_left_tc__width_256__rotation_384;
logic start__rotator_left_tc__width_256__rotation_511;
logic start__rotator_left_tc__width_256__rotation_512;

logic start__rotator_left_tc__width_512__rotation_0;
logic start__rotator_left_tc__width_512__rotation_1;
logic start__rotator_left_tc__width_512__rotation_2;
logic start__rotator_left_tc__width_512__rotation_3;
logic start__rotator_left_tc__width_512__rotation_4;
logic start__rotator_left_tc__width_512__rotation_5;
logic start__rotator_left_tc__width_512__rotation_6;
logic start__rotator_left_tc__width_512__rotation_7;
logic start__rotator_left_tc__width_512__rotation_256;
logic start__rotator_left_tc__width_512__rotation_511;
logic start__rotator_left_tc__width_512__rotation_512;
logic start__rotator_left_tc__width_512__rotation_513;
logic start__rotator_left_tc__width_512__rotation_768;
logic start__rotator_left_tc__width_512__rotation_1023;
logic start__rotator_left_tc__width_512__rotation_1024;

logic start__rotator_left_tc__width_1024__rotation_0;
logic start__rotator_left_tc__width_1024__rotation_1;
logic start__rotator_left_tc__width_1024__rotation_2;
logic start__rotator_left_tc__width_1024__rotation_3;
logic start__rotator_left_tc__width_1024__rotation_4;
logic start__rotator_left_tc__width_1024__rotation_5;
logic start__rotator_left_tc__width_1024__rotation_6;
logic start__rotator_left_tc__width_1024__rotation_7;
logic start__rotator_left_tc__width_1024__rotation_512;
logic start__rotator_left_tc__width_1024__rotation_1023;
logic start__rotator_left_tc__width_1024__rotation_1024;
logic start__rotator_left_tc__width_1024__rotation_1025;
logic start__rotator_left_tc__width_1024__rotation_1536;
logic start__rotator_left_tc__width_1024__rotation_2047;
logic start__rotator_left_tc__width_1024__rotation_2048;

rotator_left_tc #(.WIDTH(1), .ROTATION(0)) rotator_left_tc__width_1__rotation_0 (.start(start__rotator_left_tc__width_1__rotation_0));
rotator_left_tc #(.WIDTH(1), .ROTATION(1)) rotator_left_tc__width_1__rotation_1 (.start(start__rotator_left_tc__width_1__rotation_1));

rotator_left_tc #(.WIDTH(2), .ROTATION(0)) rotator_left_tc__width_2__rotation_0 (.start(start__rotator_left_tc__width_2__rotation_0));
rotator_left_tc #(.WIDTH(2), .ROTATION(1)) rotator_left_tc__width_2__rotation_1 (.start(start__rotator_left_tc__width_2__rotation_1));
rotator_left_tc #(.WIDTH(2), .ROTATION(2)) rotator_left_tc__width_2__rotation_2 (.start(start__rotator_left_tc__width_2__rotation_2));
rotator_left_tc #(.WIDTH(2), .ROTATION(3)) rotator_left_tc__width_2__rotation_3 (.start(start__rotator_left_tc__width_2__rotation_3));

rotator_left_tc #(.WIDTH(3), .ROTATION(0)) rotator_left_tc__width_3__rotation_0 (.start(start__rotator_left_tc__width_3__rotation_0));
rotator_left_tc #(.WIDTH(3), .ROTATION(1)) rotator_left_tc__width_3__rotation_1 (.start(start__rotator_left_tc__width_3__rotation_1));
rotator_left_tc #(.WIDTH(3), .ROTATION(2)) rotator_left_tc__width_3__rotation_2 (.start(start__rotator_left_tc__width_3__rotation_2));
rotator_left_tc #(.WIDTH(3), .ROTATION(3)) rotator_left_tc__width_3__rotation_3 (.start(start__rotator_left_tc__width_3__rotation_3));
rotator_left_tc #(.WIDTH(3), .ROTATION(4)) rotator_left_tc__width_3__rotation_4 (.start(start__rotator_left_tc__width_3__rotation_4));
rotator_left_tc #(.WIDTH(3), .ROTATION(5)) rotator_left_tc__width_3__rotation_5 (.start(start__rotator_left_tc__width_3__rotation_5));

rotator_left_tc #(.WIDTH(4), .ROTATION(0)) rotator_left_tc__width_4__rotation_0 (.start(start__rotator_left_tc__width_4__rotation_0));
rotator_left_tc #(.WIDTH(4), .ROTATION(1)) rotator_left_tc__width_4__rotation_1 (.start(start__rotator_left_tc__width_4__rotation_1));
rotator_left_tc #(.WIDTH(4), .ROTATION(2)) rotator_left_tc__width_4__rotation_2 (.start(start__rotator_left_tc__width_4__rotation_2));
rotator_left_tc #(.WIDTH(4), .ROTATION(3)) rotator_left_tc__width_4__rotation_3 (.start(start__rotator_left_tc__width_4__rotation_3));
rotator_left_tc #(.WIDTH(4), .ROTATION(4)) rotator_left_tc__width_4__rotation_4 (.start(start__rotator_left_tc__width_4__rotation_4));
rotator_left_tc #(.WIDTH(4), .ROTATION(5)) rotator_left_tc__width_4__rotation_5 (.start(start__rotator_left_tc__width_4__rotation_5));
rotator_left_tc #(.WIDTH(4), .ROTATION(6)) rotator_left_tc__width_4__rotation_6 (.start(start__rotator_left_tc__width_4__rotation_6));
rotator_left_tc #(.WIDTH(4), .ROTATION(7)) rotator_left_tc__width_4__rotation_7 (.start(start__rotator_left_tc__width_4__rotation_7));

rotator_left_tc #(.WIDTH(5), .ROTATION(0)) rotator_left_tc__width_5__rotation_0 (.start(start__rotator_left_tc__width_5__rotation_0));
rotator_left_tc #(.WIDTH(5), .ROTATION(1)) rotator_left_tc__width_5__rotation_1 (.start(start__rotator_left_tc__width_5__rotation_1));
rotator_left_tc #(.WIDTH(5), .ROTATION(2)) rotator_left_tc__width_5__rotation_2 (.start(start__rotator_left_tc__width_5__rotation_2));
rotator_left_tc #(.WIDTH(5), .ROTATION(3)) rotator_left_tc__width_5__rotation_3 (.start(start__rotator_left_tc__width_5__rotation_3));
rotator_left_tc #(.WIDTH(5), .ROTATION(4)) rotator_left_tc__width_5__rotation_4 (.start(start__rotator_left_tc__width_5__rotation_4));
rotator_left_tc #(.WIDTH(5), .ROTATION(5)) rotator_left_tc__width_5__rotation_5 (.start(start__rotator_left_tc__width_5__rotation_5));
rotator_left_tc #(.WIDTH(5), .ROTATION(6)) rotator_left_tc__width_5__rotation_6 (.start(start__rotator_left_tc__width_5__rotation_6));
rotator_left_tc #(.WIDTH(5), .ROTATION(7)) rotator_left_tc__width_5__rotation_7 (.start(start__rotator_left_tc__width_5__rotation_7));
rotator_left_tc #(.WIDTH(5), .ROTATION(8)) rotator_left_tc__width_5__rotation_8 (.start(start__rotator_left_tc__width_5__rotation_8));
rotator_left_tc #(.WIDTH(5), .ROTATION(9)) rotator_left_tc__width_5__rotation_9 (.start(start__rotator_left_tc__width_5__rotation_9));

rotator_left_tc #(.WIDTH(6), .ROTATION(0)) rotator_left_tc__width_6__rotation_0 (.start(start__rotator_left_tc__width_6__rotation_0));
rotator_left_tc #(.WIDTH(6), .ROTATION(1)) rotator_left_tc__width_6__rotation_1 (.start(start__rotator_left_tc__width_6__rotation_1));
rotator_left_tc #(.WIDTH(6), .ROTATION(2)) rotator_left_tc__width_6__rotation_2 (.start(start__rotator_left_tc__width_6__rotation_2));
rotator_left_tc #(.WIDTH(6), .ROTATION(3)) rotator_left_tc__width_6__rotation_3 (.start(start__rotator_left_tc__width_6__rotation_3));
rotator_left_tc #(.WIDTH(6), .ROTATION(4)) rotator_left_tc__width_6__rotation_4 (.start(start__rotator_left_tc__width_6__rotation_4));
rotator_left_tc #(.WIDTH(6), .ROTATION(5)) rotator_left_tc__width_6__rotation_5 (.start(start__rotator_left_tc__width_6__rotation_5));
rotator_left_tc #(.WIDTH(6), .ROTATION(6)) rotator_left_tc__width_6__rotation_6 (.start(start__rotator_left_tc__width_6__rotation_6));
rotator_left_tc #(.WIDTH(6), .ROTATION(7)) rotator_left_tc__width_6__rotation_7 (.start(start__rotator_left_tc__width_6__rotation_7));
rotator_left_tc #(.WIDTH(6), .ROTATION(8)) rotator_left_tc__width_6__rotation_8 (.start(start__rotator_left_tc__width_6__rotation_8));
rotator_left_tc #(.WIDTH(6), .ROTATION(9)) rotator_left_tc__width_6__rotation_9 (.start(start__rotator_left_tc__width_6__rotation_9));
rotator_left_tc #(.WIDTH(6), .ROTATION(10)) rotator_left_tc__width_6__rotation_10 (.start(start__rotator_left_tc__width_6__rotation_10));
rotator_left_tc #(.WIDTH(6), .ROTATION(11)) rotator_left_tc__width_6__rotation_11 (.start(start__rotator_left_tc__width_6__rotation_11));

rotator_left_tc #(.WIDTH(7), .ROTATION(0)) rotator_left_tc__width_7__rotation_0 (.start(start__rotator_left_tc__width_7__rotation_0));
rotator_left_tc #(.WIDTH(7), .ROTATION(1)) rotator_left_tc__width_7__rotation_1 (.start(start__rotator_left_tc__width_7__rotation_1));
rotator_left_tc #(.WIDTH(7), .ROTATION(2)) rotator_left_tc__width_7__rotation_2 (.start(start__rotator_left_tc__width_7__rotation_2));
rotator_left_tc #(.WIDTH(7), .ROTATION(3)) rotator_left_tc__width_7__rotation_3 (.start(start__rotator_left_tc__width_7__rotation_3));
rotator_left_tc #(.WIDTH(7), .ROTATION(4)) rotator_left_tc__width_7__rotation_4 (.start(start__rotator_left_tc__width_7__rotation_4));
rotator_left_tc #(.WIDTH(7), .ROTATION(5)) rotator_left_tc__width_7__rotation_5 (.start(start__rotator_left_tc__width_7__rotation_5));
rotator_left_tc #(.WIDTH(7), .ROTATION(6)) rotator_left_tc__width_7__rotation_6 (.start(start__rotator_left_tc__width_7__rotation_6));
rotator_left_tc #(.WIDTH(7), .ROTATION(7)) rotator_left_tc__width_7__rotation_7 (.start(start__rotator_left_tc__width_7__rotation_7));
rotator_left_tc #(.WIDTH(7), .ROTATION(8)) rotator_left_tc__width_7__rotation_8 (.start(start__rotator_left_tc__width_7__rotation_8));
rotator_left_tc #(.WIDTH(7), .ROTATION(9)) rotator_left_tc__width_7__rotation_9 (.start(start__rotator_left_tc__width_7__rotation_9));
rotator_left_tc #(.WIDTH(7), .ROTATION(10)) rotator_left_tc__width_7__rotation_10 (.start(start__rotator_left_tc__width_7__rotation_10));
rotator_left_tc #(.WIDTH(7), .ROTATION(11)) rotator_left_tc__width_7__rotation_11 (.start(start__rotator_left_tc__width_7__rotation_11));
rotator_left_tc #(.WIDTH(7), .ROTATION(12)) rotator_left_tc__width_7__rotation_12 (.start(start__rotator_left_tc__width_7__rotation_12));
rotator_left_tc #(.WIDTH(7), .ROTATION(13)) rotator_left_tc__width_7__rotation_13 (.start(start__rotator_left_tc__width_7__rotation_13));

rotator_left_tc #(.WIDTH(8), .ROTATION(0)) rotator_left_tc__width_8__rotation_0 (.start(start__rotator_left_tc__width_8__rotation_0));
rotator_left_tc #(.WIDTH(8), .ROTATION(1)) rotator_left_tc__width_8__rotation_1 (.start(start__rotator_left_tc__width_8__rotation_1));
rotator_left_tc #(.WIDTH(8), .ROTATION(2)) rotator_left_tc__width_8__rotation_2 (.start(start__rotator_left_tc__width_8__rotation_2));
rotator_left_tc #(.WIDTH(8), .ROTATION(3)) rotator_left_tc__width_8__rotation_3 (.start(start__rotator_left_tc__width_8__rotation_3));
rotator_left_tc #(.WIDTH(8), .ROTATION(4)) rotator_left_tc__width_8__rotation_4 (.start(start__rotator_left_tc__width_8__rotation_4));
rotator_left_tc #(.WIDTH(8), .ROTATION(5)) rotator_left_tc__width_8__rotation_5 (.start(start__rotator_left_tc__width_8__rotation_5));
rotator_left_tc #(.WIDTH(8), .ROTATION(6)) rotator_left_tc__width_8__rotation_6 (.start(start__rotator_left_tc__width_8__rotation_6));
rotator_left_tc #(.WIDTH(8), .ROTATION(7)) rotator_left_tc__width_8__rotation_7 (.start(start__rotator_left_tc__width_8__rotation_7));
rotator_left_tc #(.WIDTH(8), .ROTATION(8)) rotator_left_tc__width_8__rotation_8 (.start(start__rotator_left_tc__width_8__rotation_8));
rotator_left_tc #(.WIDTH(8), .ROTATION(9)) rotator_left_tc__width_8__rotation_9 (.start(start__rotator_left_tc__width_8__rotation_9));
rotator_left_tc #(.WIDTH(8), .ROTATION(10)) rotator_left_tc__width_8__rotation_10 (.start(start__rotator_left_tc__width_8__rotation_10));
rotator_left_tc #(.WIDTH(8), .ROTATION(11)) rotator_left_tc__width_8__rotation_11 (.start(start__rotator_left_tc__width_8__rotation_11));
rotator_left_tc #(.WIDTH(8), .ROTATION(12)) rotator_left_tc__width_8__rotation_12 (.start(start__rotator_left_tc__width_8__rotation_12));
rotator_left_tc #(.WIDTH(8), .ROTATION(13)) rotator_left_tc__width_8__rotation_13 (.start(start__rotator_left_tc__width_8__rotation_13));
rotator_left_tc #(.WIDTH(8), .ROTATION(14)) rotator_left_tc__width_8__rotation_14 (.start(start__rotator_left_tc__width_8__rotation_14));
rotator_left_tc #(.WIDTH(8), .ROTATION(15)) rotator_left_tc__width_8__rotation_15 (.start(start__rotator_left_tc__width_8__rotation_15));

rotator_left_tc #(.WIDTH(9), .ROTATION(0)) rotator_left_tc__width_9__rotation_0 (.start(start__rotator_left_tc__width_9__rotation_0));
rotator_left_tc #(.WIDTH(9), .ROTATION(1)) rotator_left_tc__width_9__rotation_1 (.start(start__rotator_left_tc__width_9__rotation_1));
rotator_left_tc #(.WIDTH(9), .ROTATION(2)) rotator_left_tc__width_9__rotation_2 (.start(start__rotator_left_tc__width_9__rotation_2));
rotator_left_tc #(.WIDTH(9), .ROTATION(3)) rotator_left_tc__width_9__rotation_3 (.start(start__rotator_left_tc__width_9__rotation_3));
rotator_left_tc #(.WIDTH(9), .ROTATION(4)) rotator_left_tc__width_9__rotation_4 (.start(start__rotator_left_tc__width_9__rotation_4));
rotator_left_tc #(.WIDTH(9), .ROTATION(5)) rotator_left_tc__width_9__rotation_5 (.start(start__rotator_left_tc__width_9__rotation_5));
rotator_left_tc #(.WIDTH(9), .ROTATION(6)) rotator_left_tc__width_9__rotation_6 (.start(start__rotator_left_tc__width_9__rotation_6));
rotator_left_tc #(.WIDTH(9), .ROTATION(7)) rotator_left_tc__width_9__rotation_7 (.start(start__rotator_left_tc__width_9__rotation_7));
rotator_left_tc #(.WIDTH(9), .ROTATION(8)) rotator_left_tc__width_9__rotation_8 (.start(start__rotator_left_tc__width_9__rotation_8));
rotator_left_tc #(.WIDTH(9), .ROTATION(9)) rotator_left_tc__width_9__rotation_9 (.start(start__rotator_left_tc__width_9__rotation_9));
rotator_left_tc #(.WIDTH(9), .ROTATION(10)) rotator_left_tc__width_9__rotation_10 (.start(start__rotator_left_tc__width_9__rotation_10));
rotator_left_tc #(.WIDTH(9), .ROTATION(11)) rotator_left_tc__width_9__rotation_11 (.start(start__rotator_left_tc__width_9__rotation_11));
rotator_left_tc #(.WIDTH(9), .ROTATION(12)) rotator_left_tc__width_9__rotation_12 (.start(start__rotator_left_tc__width_9__rotation_12));
rotator_left_tc #(.WIDTH(9), .ROTATION(13)) rotator_left_tc__width_9__rotation_13 (.start(start__rotator_left_tc__width_9__rotation_13));
rotator_left_tc #(.WIDTH(9), .ROTATION(14)) rotator_left_tc__width_9__rotation_14 (.start(start__rotator_left_tc__width_9__rotation_14));
rotator_left_tc #(.WIDTH(9), .ROTATION(15)) rotator_left_tc__width_9__rotation_15 (.start(start__rotator_left_tc__width_9__rotation_15));
rotator_left_tc #(.WIDTH(9), .ROTATION(16)) rotator_left_tc__width_9__rotation_16 (.start(start__rotator_left_tc__width_9__rotation_16));
rotator_left_tc #(.WIDTH(9), .ROTATION(17)) rotator_left_tc__width_9__rotation_17 (.start(start__rotator_left_tc__width_9__rotation_17));

rotator_left_tc #(.WIDTH(10), .ROTATION(0)) rotator_left_tc__width_10__rotation_0 (.start(start__rotator_left_tc__width_10__rotation_0));
rotator_left_tc #(.WIDTH(10), .ROTATION(1)) rotator_left_tc__width_10__rotation_1 (.start(start__rotator_left_tc__width_10__rotation_1));
rotator_left_tc #(.WIDTH(10), .ROTATION(2)) rotator_left_tc__width_10__rotation_2 (.start(start__rotator_left_tc__width_10__rotation_2));
rotator_left_tc #(.WIDTH(10), .ROTATION(3)) rotator_left_tc__width_10__rotation_3 (.start(start__rotator_left_tc__width_10__rotation_3));
rotator_left_tc #(.WIDTH(10), .ROTATION(4)) rotator_left_tc__width_10__rotation_4 (.start(start__rotator_left_tc__width_10__rotation_4));
rotator_left_tc #(.WIDTH(10), .ROTATION(5)) rotator_left_tc__width_10__rotation_5 (.start(start__rotator_left_tc__width_10__rotation_5));
rotator_left_tc #(.WIDTH(10), .ROTATION(6)) rotator_left_tc__width_10__rotation_6 (.start(start__rotator_left_tc__width_10__rotation_6));
rotator_left_tc #(.WIDTH(10), .ROTATION(7)) rotator_left_tc__width_10__rotation_7 (.start(start__rotator_left_tc__width_10__rotation_7));
rotator_left_tc #(.WIDTH(10), .ROTATION(8)) rotator_left_tc__width_10__rotation_8 (.start(start__rotator_left_tc__width_10__rotation_8));
rotator_left_tc #(.WIDTH(10), .ROTATION(9)) rotator_left_tc__width_10__rotation_9 (.start(start__rotator_left_tc__width_10__rotation_9));
rotator_left_tc #(.WIDTH(10), .ROTATION(10)) rotator_left_tc__width_10__rotation_10 (.start(start__rotator_left_tc__width_10__rotation_10));
rotator_left_tc #(.WIDTH(10), .ROTATION(11)) rotator_left_tc__width_10__rotation_11 (.start(start__rotator_left_tc__width_10__rotation_11));
rotator_left_tc #(.WIDTH(10), .ROTATION(12)) rotator_left_tc__width_10__rotation_12 (.start(start__rotator_left_tc__width_10__rotation_12));
rotator_left_tc #(.WIDTH(10), .ROTATION(13)) rotator_left_tc__width_10__rotation_13 (.start(start__rotator_left_tc__width_10__rotation_13));
rotator_left_tc #(.WIDTH(10), .ROTATION(14)) rotator_left_tc__width_10__rotation_14 (.start(start__rotator_left_tc__width_10__rotation_14));
rotator_left_tc #(.WIDTH(10), .ROTATION(15)) rotator_left_tc__width_10__rotation_15 (.start(start__rotator_left_tc__width_10__rotation_15));
rotator_left_tc #(.WIDTH(10), .ROTATION(16)) rotator_left_tc__width_10__rotation_16 (.start(start__rotator_left_tc__width_10__rotation_16));
rotator_left_tc #(.WIDTH(10), .ROTATION(17)) rotator_left_tc__width_10__rotation_17 (.start(start__rotator_left_tc__width_10__rotation_17));
rotator_left_tc #(.WIDTH(10), .ROTATION(18)) rotator_left_tc__width_10__rotation_18 (.start(start__rotator_left_tc__width_10__rotation_18));
rotator_left_tc #(.WIDTH(10), .ROTATION(19)) rotator_left_tc__width_10__rotation_19 (.start(start__rotator_left_tc__width_10__rotation_19));

rotator_left_tc #(.WIDTH(11), .ROTATION(0)) rotator_left_tc__width_11__rotation_0 (.start(start__rotator_left_tc__width_11__rotation_0));
rotator_left_tc #(.WIDTH(11), .ROTATION(1)) rotator_left_tc__width_11__rotation_1 (.start(start__rotator_left_tc__width_11__rotation_1));
rotator_left_tc #(.WIDTH(11), .ROTATION(2)) rotator_left_tc__width_11__rotation_2 (.start(start__rotator_left_tc__width_11__rotation_2));
rotator_left_tc #(.WIDTH(11), .ROTATION(3)) rotator_left_tc__width_11__rotation_3 (.start(start__rotator_left_tc__width_11__rotation_3));
rotator_left_tc #(.WIDTH(11), .ROTATION(4)) rotator_left_tc__width_11__rotation_4 (.start(start__rotator_left_tc__width_11__rotation_4));
rotator_left_tc #(.WIDTH(11), .ROTATION(5)) rotator_left_tc__width_11__rotation_5 (.start(start__rotator_left_tc__width_11__rotation_5));
rotator_left_tc #(.WIDTH(11), .ROTATION(6)) rotator_left_tc__width_11__rotation_6 (.start(start__rotator_left_tc__width_11__rotation_6));
rotator_left_tc #(.WIDTH(11), .ROTATION(7)) rotator_left_tc__width_11__rotation_7 (.start(start__rotator_left_tc__width_11__rotation_7));
rotator_left_tc #(.WIDTH(11), .ROTATION(8)) rotator_left_tc__width_11__rotation_8 (.start(start__rotator_left_tc__width_11__rotation_8));
rotator_left_tc #(.WIDTH(11), .ROTATION(9)) rotator_left_tc__width_11__rotation_9 (.start(start__rotator_left_tc__width_11__rotation_9));
rotator_left_tc #(.WIDTH(11), .ROTATION(10)) rotator_left_tc__width_11__rotation_10 (.start(start__rotator_left_tc__width_11__rotation_10));
rotator_left_tc #(.WIDTH(11), .ROTATION(11)) rotator_left_tc__width_11__rotation_11 (.start(start__rotator_left_tc__width_11__rotation_11));
rotator_left_tc #(.WIDTH(11), .ROTATION(12)) rotator_left_tc__width_11__rotation_12 (.start(start__rotator_left_tc__width_11__rotation_12));
rotator_left_tc #(.WIDTH(11), .ROTATION(13)) rotator_left_tc__width_11__rotation_13 (.start(start__rotator_left_tc__width_11__rotation_13));
rotator_left_tc #(.WIDTH(11), .ROTATION(14)) rotator_left_tc__width_11__rotation_14 (.start(start__rotator_left_tc__width_11__rotation_14));
rotator_left_tc #(.WIDTH(11), .ROTATION(15)) rotator_left_tc__width_11__rotation_15 (.start(start__rotator_left_tc__width_11__rotation_15));
rotator_left_tc #(.WIDTH(11), .ROTATION(16)) rotator_left_tc__width_11__rotation_16 (.start(start__rotator_left_tc__width_11__rotation_16));
rotator_left_tc #(.WIDTH(11), .ROTATION(17)) rotator_left_tc__width_11__rotation_17 (.start(start__rotator_left_tc__width_11__rotation_17));
rotator_left_tc #(.WIDTH(11), .ROTATION(18)) rotator_left_tc__width_11__rotation_18 (.start(start__rotator_left_tc__width_11__rotation_18));
rotator_left_tc #(.WIDTH(11), .ROTATION(19)) rotator_left_tc__width_11__rotation_19 (.start(start__rotator_left_tc__width_11__rotation_19));
rotator_left_tc #(.WIDTH(11), .ROTATION(20)) rotator_left_tc__width_11__rotation_20 (.start(start__rotator_left_tc__width_11__rotation_20));
rotator_left_tc #(.WIDTH(11), .ROTATION(21)) rotator_left_tc__width_11__rotation_21 (.start(start__rotator_left_tc__width_11__rotation_21));

rotator_left_tc #(.WIDTH(12), .ROTATION(0)) rotator_left_tc__width_12__rotation_0 (.start(start__rotator_left_tc__width_12__rotation_0));
rotator_left_tc #(.WIDTH(12), .ROTATION(1)) rotator_left_tc__width_12__rotation_1 (.start(start__rotator_left_tc__width_12__rotation_1));
rotator_left_tc #(.WIDTH(12), .ROTATION(2)) rotator_left_tc__width_12__rotation_2 (.start(start__rotator_left_tc__width_12__rotation_2));
rotator_left_tc #(.WIDTH(12), .ROTATION(3)) rotator_left_tc__width_12__rotation_3 (.start(start__rotator_left_tc__width_12__rotation_3));
rotator_left_tc #(.WIDTH(12), .ROTATION(4)) rotator_left_tc__width_12__rotation_4 (.start(start__rotator_left_tc__width_12__rotation_4));
rotator_left_tc #(.WIDTH(12), .ROTATION(5)) rotator_left_tc__width_12__rotation_5 (.start(start__rotator_left_tc__width_12__rotation_5));
rotator_left_tc #(.WIDTH(12), .ROTATION(6)) rotator_left_tc__width_12__rotation_6 (.start(start__rotator_left_tc__width_12__rotation_6));
rotator_left_tc #(.WIDTH(12), .ROTATION(7)) rotator_left_tc__width_12__rotation_7 (.start(start__rotator_left_tc__width_12__rotation_7));
rotator_left_tc #(.WIDTH(12), .ROTATION(8)) rotator_left_tc__width_12__rotation_8 (.start(start__rotator_left_tc__width_12__rotation_8));
rotator_left_tc #(.WIDTH(12), .ROTATION(9)) rotator_left_tc__width_12__rotation_9 (.start(start__rotator_left_tc__width_12__rotation_9));
rotator_left_tc #(.WIDTH(12), .ROTATION(10)) rotator_left_tc__width_12__rotation_10 (.start(start__rotator_left_tc__width_12__rotation_10));
rotator_left_tc #(.WIDTH(12), .ROTATION(11)) rotator_left_tc__width_12__rotation_11 (.start(start__rotator_left_tc__width_12__rotation_11));
rotator_left_tc #(.WIDTH(12), .ROTATION(12)) rotator_left_tc__width_12__rotation_12 (.start(start__rotator_left_tc__width_12__rotation_12));
rotator_left_tc #(.WIDTH(12), .ROTATION(13)) rotator_left_tc__width_12__rotation_13 (.start(start__rotator_left_tc__width_12__rotation_13));
rotator_left_tc #(.WIDTH(12), .ROTATION(14)) rotator_left_tc__width_12__rotation_14 (.start(start__rotator_left_tc__width_12__rotation_14));
rotator_left_tc #(.WIDTH(12), .ROTATION(15)) rotator_left_tc__width_12__rotation_15 (.start(start__rotator_left_tc__width_12__rotation_15));
rotator_left_tc #(.WIDTH(12), .ROTATION(16)) rotator_left_tc__width_12__rotation_16 (.start(start__rotator_left_tc__width_12__rotation_16));
rotator_left_tc #(.WIDTH(12), .ROTATION(17)) rotator_left_tc__width_12__rotation_17 (.start(start__rotator_left_tc__width_12__rotation_17));
rotator_left_tc #(.WIDTH(12), .ROTATION(18)) rotator_left_tc__width_12__rotation_18 (.start(start__rotator_left_tc__width_12__rotation_18));
rotator_left_tc #(.WIDTH(12), .ROTATION(19)) rotator_left_tc__width_12__rotation_19 (.start(start__rotator_left_tc__width_12__rotation_19));
rotator_left_tc #(.WIDTH(12), .ROTATION(20)) rotator_left_tc__width_12__rotation_20 (.start(start__rotator_left_tc__width_12__rotation_20));
rotator_left_tc #(.WIDTH(12), .ROTATION(21)) rotator_left_tc__width_12__rotation_21 (.start(start__rotator_left_tc__width_12__rotation_21));
rotator_left_tc #(.WIDTH(12), .ROTATION(22)) rotator_left_tc__width_12__rotation_22 (.start(start__rotator_left_tc__width_12__rotation_22));
rotator_left_tc #(.WIDTH(12), .ROTATION(23)) rotator_left_tc__width_12__rotation_23 (.start(start__rotator_left_tc__width_12__rotation_23));

rotator_left_tc #(.WIDTH(16), .ROTATION(0)) rotator_left_tc__width_16__rotation_0 (.start(start__rotator_left_tc__width_16__rotation_0));
rotator_left_tc #(.WIDTH(16), .ROTATION(1)) rotator_left_tc__width_16__rotation_1 (.start(start__rotator_left_tc__width_16__rotation_1));
rotator_left_tc #(.WIDTH(16), .ROTATION(2)) rotator_left_tc__width_16__rotation_2 (.start(start__rotator_left_tc__width_16__rotation_2));
rotator_left_tc #(.WIDTH(16), .ROTATION(3)) rotator_left_tc__width_16__rotation_3 (.start(start__rotator_left_tc__width_16__rotation_3));
rotator_left_tc #(.WIDTH(16), .ROTATION(4)) rotator_left_tc__width_16__rotation_4 (.start(start__rotator_left_tc__width_16__rotation_4));
rotator_left_tc #(.WIDTH(16), .ROTATION(5)) rotator_left_tc__width_16__rotation_5 (.start(start__rotator_left_tc__width_16__rotation_5));
rotator_left_tc #(.WIDTH(16), .ROTATION(6)) rotator_left_tc__width_16__rotation_6 (.start(start__rotator_left_tc__width_16__rotation_6));
rotator_left_tc #(.WIDTH(16), .ROTATION(7)) rotator_left_tc__width_16__rotation_7 (.start(start__rotator_left_tc__width_16__rotation_7));
rotator_left_tc #(.WIDTH(16), .ROTATION(8)) rotator_left_tc__width_16__rotation_8 (.start(start__rotator_left_tc__width_16__rotation_8));
rotator_left_tc #(.WIDTH(16), .ROTATION(15)) rotator_left_tc__width_16__rotation_15 (.start(start__rotator_left_tc__width_16__rotation_15));
rotator_left_tc #(.WIDTH(16), .ROTATION(16)) rotator_left_tc__width_16__rotation_16 (.start(start__rotator_left_tc__width_16__rotation_16));
rotator_left_tc #(.WIDTH(16), .ROTATION(17)) rotator_left_tc__width_16__rotation_17 (.start(start__rotator_left_tc__width_16__rotation_17));
rotator_left_tc #(.WIDTH(16), .ROTATION(24)) rotator_left_tc__width_16__rotation_24 (.start(start__rotator_left_tc__width_16__rotation_24));
rotator_left_tc #(.WIDTH(16), .ROTATION(31)) rotator_left_tc__width_16__rotation_31 (.start(start__rotator_left_tc__width_16__rotation_31));
rotator_left_tc #(.WIDTH(16), .ROTATION(32)) rotator_left_tc__width_16__rotation_32 (.start(start__rotator_left_tc__width_16__rotation_32));

rotator_left_tc #(.WIDTH(24), .ROTATION(0)) rotator_left_tc__width_24__rotation_0 (.start(start__rotator_left_tc__width_24__rotation_0));
rotator_left_tc #(.WIDTH(24), .ROTATION(1)) rotator_left_tc__width_24__rotation_1 (.start(start__rotator_left_tc__width_24__rotation_1));
rotator_left_tc #(.WIDTH(24), .ROTATION(2)) rotator_left_tc__width_24__rotation_2 (.start(start__rotator_left_tc__width_24__rotation_2));
rotator_left_tc #(.WIDTH(24), .ROTATION(3)) rotator_left_tc__width_24__rotation_3 (.start(start__rotator_left_tc__width_24__rotation_3));
rotator_left_tc #(.WIDTH(24), .ROTATION(4)) rotator_left_tc__width_24__rotation_4 (.start(start__rotator_left_tc__width_24__rotation_4));
rotator_left_tc #(.WIDTH(24), .ROTATION(5)) rotator_left_tc__width_24__rotation_5 (.start(start__rotator_left_tc__width_24__rotation_5));
rotator_left_tc #(.WIDTH(24), .ROTATION(6)) rotator_left_tc__width_24__rotation_6 (.start(start__rotator_left_tc__width_24__rotation_6));
rotator_left_tc #(.WIDTH(24), .ROTATION(7)) rotator_left_tc__width_24__rotation_7 (.start(start__rotator_left_tc__width_24__rotation_7));
rotator_left_tc #(.WIDTH(24), .ROTATION(12)) rotator_left_tc__width_24__rotation_12 (.start(start__rotator_left_tc__width_24__rotation_12));
rotator_left_tc #(.WIDTH(24), .ROTATION(23)) rotator_left_tc__width_24__rotation_23 (.start(start__rotator_left_tc__width_24__rotation_23));
rotator_left_tc #(.WIDTH(24), .ROTATION(24)) rotator_left_tc__width_24__rotation_24 (.start(start__rotator_left_tc__width_24__rotation_24));
rotator_left_tc #(.WIDTH(24), .ROTATION(25)) rotator_left_tc__width_24__rotation_25 (.start(start__rotator_left_tc__width_24__rotation_25));
rotator_left_tc #(.WIDTH(24), .ROTATION(36)) rotator_left_tc__width_24__rotation_36 (.start(start__rotator_left_tc__width_24__rotation_36));
rotator_left_tc #(.WIDTH(24), .ROTATION(47)) rotator_left_tc__width_24__rotation_47 (.start(start__rotator_left_tc__width_24__rotation_47));
rotator_left_tc #(.WIDTH(24), .ROTATION(48)) rotator_left_tc__width_24__rotation_48 (.start(start__rotator_left_tc__width_24__rotation_48));

rotator_left_tc #(.WIDTH(32), .ROTATION(0)) rotator_left_tc__width_32__rotation_0 (.start(start__rotator_left_tc__width_32__rotation_0));
rotator_left_tc #(.WIDTH(32), .ROTATION(1)) rotator_left_tc__width_32__rotation_1 (.start(start__rotator_left_tc__width_32__rotation_1));
rotator_left_tc #(.WIDTH(32), .ROTATION(2)) rotator_left_tc__width_32__rotation_2 (.start(start__rotator_left_tc__width_32__rotation_2));
rotator_left_tc #(.WIDTH(32), .ROTATION(3)) rotator_left_tc__width_32__rotation_3 (.start(start__rotator_left_tc__width_32__rotation_3));
rotator_left_tc #(.WIDTH(32), .ROTATION(4)) rotator_left_tc__width_32__rotation_4 (.start(start__rotator_left_tc__width_32__rotation_4));
rotator_left_tc #(.WIDTH(32), .ROTATION(5)) rotator_left_tc__width_32__rotation_5 (.start(start__rotator_left_tc__width_32__rotation_5));
rotator_left_tc #(.WIDTH(32), .ROTATION(6)) rotator_left_tc__width_32__rotation_6 (.start(start__rotator_left_tc__width_32__rotation_6));
rotator_left_tc #(.WIDTH(32), .ROTATION(7)) rotator_left_tc__width_32__rotation_7 (.start(start__rotator_left_tc__width_32__rotation_7));
rotator_left_tc #(.WIDTH(32), .ROTATION(16)) rotator_left_tc__width_32__rotation_16 (.start(start__rotator_left_tc__width_32__rotation_16));
rotator_left_tc #(.WIDTH(32), .ROTATION(31)) rotator_left_tc__width_32__rotation_31 (.start(start__rotator_left_tc__width_32__rotation_31));
rotator_left_tc #(.WIDTH(32), .ROTATION(32)) rotator_left_tc__width_32__rotation_32 (.start(start__rotator_left_tc__width_32__rotation_32));
rotator_left_tc #(.WIDTH(32), .ROTATION(33)) rotator_left_tc__width_32__rotation_33 (.start(start__rotator_left_tc__width_32__rotation_33));
rotator_left_tc #(.WIDTH(32), .ROTATION(48)) rotator_left_tc__width_32__rotation_48 (.start(start__rotator_left_tc__width_32__rotation_48));
rotator_left_tc #(.WIDTH(32), .ROTATION(63)) rotator_left_tc__width_32__rotation_63 (.start(start__rotator_left_tc__width_32__rotation_63));
rotator_left_tc #(.WIDTH(32), .ROTATION(64)) rotator_left_tc__width_32__rotation_64 (.start(start__rotator_left_tc__width_32__rotation_64));

rotator_left_tc #(.WIDTH(48), .ROTATION(0)) rotator_left_tc__width_48__rotation_0 (.start(start__rotator_left_tc__width_48__rotation_0));
rotator_left_tc #(.WIDTH(48), .ROTATION(1)) rotator_left_tc__width_48__rotation_1 (.start(start__rotator_left_tc__width_48__rotation_1));
rotator_left_tc #(.WIDTH(48), .ROTATION(2)) rotator_left_tc__width_48__rotation_2 (.start(start__rotator_left_tc__width_48__rotation_2));
rotator_left_tc #(.WIDTH(48), .ROTATION(3)) rotator_left_tc__width_48__rotation_3 (.start(start__rotator_left_tc__width_48__rotation_3));
rotator_left_tc #(.WIDTH(48), .ROTATION(4)) rotator_left_tc__width_48__rotation_4 (.start(start__rotator_left_tc__width_48__rotation_4));
rotator_left_tc #(.WIDTH(48), .ROTATION(5)) rotator_left_tc__width_48__rotation_5 (.start(start__rotator_left_tc__width_48__rotation_5));
rotator_left_tc #(.WIDTH(48), .ROTATION(6)) rotator_left_tc__width_48__rotation_6 (.start(start__rotator_left_tc__width_48__rotation_6));
rotator_left_tc #(.WIDTH(48), .ROTATION(7)) rotator_left_tc__width_48__rotation_7 (.start(start__rotator_left_tc__width_48__rotation_7));
rotator_left_tc #(.WIDTH(48), .ROTATION(24)) rotator_left_tc__width_48__rotation_24 (.start(start__rotator_left_tc__width_48__rotation_24));
rotator_left_tc #(.WIDTH(48), .ROTATION(47)) rotator_left_tc__width_48__rotation_47 (.start(start__rotator_left_tc__width_48__rotation_47));
rotator_left_tc #(.WIDTH(48), .ROTATION(48)) rotator_left_tc__width_48__rotation_48 (.start(start__rotator_left_tc__width_48__rotation_48));
rotator_left_tc #(.WIDTH(48), .ROTATION(49)) rotator_left_tc__width_48__rotation_49 (.start(start__rotator_left_tc__width_48__rotation_49));
rotator_left_tc #(.WIDTH(48), .ROTATION(72)) rotator_left_tc__width_48__rotation_72 (.start(start__rotator_left_tc__width_48__rotation_72));
rotator_left_tc #(.WIDTH(48), .ROTATION(95)) rotator_left_tc__width_48__rotation_95 (.start(start__rotator_left_tc__width_48__rotation_95));
rotator_left_tc #(.WIDTH(48), .ROTATION(96)) rotator_left_tc__width_48__rotation_96 (.start(start__rotator_left_tc__width_48__rotation_96));

rotator_left_tc #(.WIDTH(64), .ROTATION(0)) rotator_left_tc__width_64__rotation_0 (.start(start__rotator_left_tc__width_64__rotation_0));
rotator_left_tc #(.WIDTH(64), .ROTATION(1)) rotator_left_tc__width_64__rotation_1 (.start(start__rotator_left_tc__width_64__rotation_1));
rotator_left_tc #(.WIDTH(64), .ROTATION(2)) rotator_left_tc__width_64__rotation_2 (.start(start__rotator_left_tc__width_64__rotation_2));
rotator_left_tc #(.WIDTH(64), .ROTATION(3)) rotator_left_tc__width_64__rotation_3 (.start(start__rotator_left_tc__width_64__rotation_3));
rotator_left_tc #(.WIDTH(64), .ROTATION(4)) rotator_left_tc__width_64__rotation_4 (.start(start__rotator_left_tc__width_64__rotation_4));
rotator_left_tc #(.WIDTH(64), .ROTATION(5)) rotator_left_tc__width_64__rotation_5 (.start(start__rotator_left_tc__width_64__rotation_5));
rotator_left_tc #(.WIDTH(64), .ROTATION(6)) rotator_left_tc__width_64__rotation_6 (.start(start__rotator_left_tc__width_64__rotation_6));
rotator_left_tc #(.WIDTH(64), .ROTATION(7)) rotator_left_tc__width_64__rotation_7 (.start(start__rotator_left_tc__width_64__rotation_7));
rotator_left_tc #(.WIDTH(64), .ROTATION(32)) rotator_left_tc__width_64__rotation_32 (.start(start__rotator_left_tc__width_64__rotation_32));
rotator_left_tc #(.WIDTH(64), .ROTATION(63)) rotator_left_tc__width_64__rotation_63 (.start(start__rotator_left_tc__width_64__rotation_63));
rotator_left_tc #(.WIDTH(64), .ROTATION(64)) rotator_left_tc__width_64__rotation_64 (.start(start__rotator_left_tc__width_64__rotation_64));
rotator_left_tc #(.WIDTH(64), .ROTATION(65)) rotator_left_tc__width_64__rotation_65 (.start(start__rotator_left_tc__width_64__rotation_65));
rotator_left_tc #(.WIDTH(64), .ROTATION(96)) rotator_left_tc__width_64__rotation_96 (.start(start__rotator_left_tc__width_64__rotation_96));
rotator_left_tc #(.WIDTH(64), .ROTATION(127)) rotator_left_tc__width_64__rotation_127 (.start(start__rotator_left_tc__width_64__rotation_127));
rotator_left_tc #(.WIDTH(64), .ROTATION(128)) rotator_left_tc__width_64__rotation_128 (.start(start__rotator_left_tc__width_64__rotation_128));

rotator_left_tc #(.WIDTH(128), .ROTATION(0)) rotator_left_tc__width_128__rotation_0 (.start(start__rotator_left_tc__width_128__rotation_0));
rotator_left_tc #(.WIDTH(128), .ROTATION(1)) rotator_left_tc__width_128__rotation_1 (.start(start__rotator_left_tc__width_128__rotation_1));
rotator_left_tc #(.WIDTH(128), .ROTATION(2)) rotator_left_tc__width_128__rotation_2 (.start(start__rotator_left_tc__width_128__rotation_2));
rotator_left_tc #(.WIDTH(128), .ROTATION(3)) rotator_left_tc__width_128__rotation_3 (.start(start__rotator_left_tc__width_128__rotation_3));
rotator_left_tc #(.WIDTH(128), .ROTATION(4)) rotator_left_tc__width_128__rotation_4 (.start(start__rotator_left_tc__width_128__rotation_4));
rotator_left_tc #(.WIDTH(128), .ROTATION(5)) rotator_left_tc__width_128__rotation_5 (.start(start__rotator_left_tc__width_128__rotation_5));
rotator_left_tc #(.WIDTH(128), .ROTATION(6)) rotator_left_tc__width_128__rotation_6 (.start(start__rotator_left_tc__width_128__rotation_6));
rotator_left_tc #(.WIDTH(128), .ROTATION(7)) rotator_left_tc__width_128__rotation_7 (.start(start__rotator_left_tc__width_128__rotation_7));
rotator_left_tc #(.WIDTH(128), .ROTATION(64)) rotator_left_tc__width_128__rotation_64 (.start(start__rotator_left_tc__width_128__rotation_64));
rotator_left_tc #(.WIDTH(128), .ROTATION(127)) rotator_left_tc__width_128__rotation_127 (.start(start__rotator_left_tc__width_128__rotation_127));
rotator_left_tc #(.WIDTH(128), .ROTATION(128)) rotator_left_tc__width_128__rotation_128 (.start(start__rotator_left_tc__width_128__rotation_128));
rotator_left_tc #(.WIDTH(128), .ROTATION(129)) rotator_left_tc__width_128__rotation_129 (.start(start__rotator_left_tc__width_128__rotation_129));
rotator_left_tc #(.WIDTH(128), .ROTATION(192)) rotator_left_tc__width_128__rotation_192 (.start(start__rotator_left_tc__width_128__rotation_192));
rotator_left_tc #(.WIDTH(128), .ROTATION(255)) rotator_left_tc__width_128__rotation_255 (.start(start__rotator_left_tc__width_128__rotation_255));
rotator_left_tc #(.WIDTH(128), .ROTATION(256)) rotator_left_tc__width_128__rotation_256 (.start(start__rotator_left_tc__width_128__rotation_256));

rotator_left_tc #(.WIDTH(256), .ROTATION(0)) rotator_left_tc__width_256__rotation_0 (.start(start__rotator_left_tc__width_256__rotation_0));
rotator_left_tc #(.WIDTH(256), .ROTATION(1)) rotator_left_tc__width_256__rotation_1 (.start(start__rotator_left_tc__width_256__rotation_1));
rotator_left_tc #(.WIDTH(256), .ROTATION(2)) rotator_left_tc__width_256__rotation_2 (.start(start__rotator_left_tc__width_256__rotation_2));
rotator_left_tc #(.WIDTH(256), .ROTATION(3)) rotator_left_tc__width_256__rotation_3 (.start(start__rotator_left_tc__width_256__rotation_3));
rotator_left_tc #(.WIDTH(256), .ROTATION(4)) rotator_left_tc__width_256__rotation_4 (.start(start__rotator_left_tc__width_256__rotation_4));
rotator_left_tc #(.WIDTH(256), .ROTATION(5)) rotator_left_tc__width_256__rotation_5 (.start(start__rotator_left_tc__width_256__rotation_5));
rotator_left_tc #(.WIDTH(256), .ROTATION(6)) rotator_left_tc__width_256__rotation_6 (.start(start__rotator_left_tc__width_256__rotation_6));
rotator_left_tc #(.WIDTH(256), .ROTATION(7)) rotator_left_tc__width_256__rotation_7 (.start(start__rotator_left_tc__width_256__rotation_7));
rotator_left_tc #(.WIDTH(256), .ROTATION(128)) rotator_left_tc__width_256__rotation_128 (.start(start__rotator_left_tc__width_256__rotation_128));
rotator_left_tc #(.WIDTH(256), .ROTATION(255)) rotator_left_tc__width_256__rotation_255 (.start(start__rotator_left_tc__width_256__rotation_255));
rotator_left_tc #(.WIDTH(256), .ROTATION(256)) rotator_left_tc__width_256__rotation_256 (.start(start__rotator_left_tc__width_256__rotation_256));
rotator_left_tc #(.WIDTH(256), .ROTATION(257)) rotator_left_tc__width_256__rotation_257 (.start(start__rotator_left_tc__width_256__rotation_257));
rotator_left_tc #(.WIDTH(256), .ROTATION(384)) rotator_left_tc__width_256__rotation_384 (.start(start__rotator_left_tc__width_256__rotation_384));
rotator_left_tc #(.WIDTH(256), .ROTATION(511)) rotator_left_tc__width_256__rotation_511 (.start(start__rotator_left_tc__width_256__rotation_511));
rotator_left_tc #(.WIDTH(256), .ROTATION(512)) rotator_left_tc__width_256__rotation_512 (.start(start__rotator_left_tc__width_256__rotation_512));

rotator_left_tc #(.WIDTH(512), .ROTATION(0)) rotator_left_tc__width_512__rotation_0 (.start(start__rotator_left_tc__width_512__rotation_0));
rotator_left_tc #(.WIDTH(512), .ROTATION(1)) rotator_left_tc__width_512__rotation_1 (.start(start__rotator_left_tc__width_512__rotation_1));
rotator_left_tc #(.WIDTH(512), .ROTATION(2)) rotator_left_tc__width_512__rotation_2 (.start(start__rotator_left_tc__width_512__rotation_2));
rotator_left_tc #(.WIDTH(512), .ROTATION(3)) rotator_left_tc__width_512__rotation_3 (.start(start__rotator_left_tc__width_512__rotation_3));
rotator_left_tc #(.WIDTH(512), .ROTATION(4)) rotator_left_tc__width_512__rotation_4 (.start(start__rotator_left_tc__width_512__rotation_4));
rotator_left_tc #(.WIDTH(512), .ROTATION(5)) rotator_left_tc__width_512__rotation_5 (.start(start__rotator_left_tc__width_512__rotation_5));
rotator_left_tc #(.WIDTH(512), .ROTATION(6)) rotator_left_tc__width_512__rotation_6 (.start(start__rotator_left_tc__width_512__rotation_6));
rotator_left_tc #(.WIDTH(512), .ROTATION(7)) rotator_left_tc__width_512__rotation_7 (.start(start__rotator_left_tc__width_512__rotation_7));
rotator_left_tc #(.WIDTH(512), .ROTATION(256)) rotator_left_tc__width_512__rotation_256 (.start(start__rotator_left_tc__width_512__rotation_256));
rotator_left_tc #(.WIDTH(512), .ROTATION(511)) rotator_left_tc__width_512__rotation_511 (.start(start__rotator_left_tc__width_512__rotation_511));
rotator_left_tc #(.WIDTH(512), .ROTATION(512)) rotator_left_tc__width_512__rotation_512 (.start(start__rotator_left_tc__width_512__rotation_512));
rotator_left_tc #(.WIDTH(512), .ROTATION(513)) rotator_left_tc__width_512__rotation_513 (.start(start__rotator_left_tc__width_512__rotation_513));
rotator_left_tc #(.WIDTH(512), .ROTATION(768)) rotator_left_tc__width_512__rotation_768 (.start(start__rotator_left_tc__width_512__rotation_768));
rotator_left_tc #(.WIDTH(512), .ROTATION(1023)) rotator_left_tc__width_512__rotation_1023 (.start(start__rotator_left_tc__width_512__rotation_1023));
rotator_left_tc #(.WIDTH(512), .ROTATION(1024)) rotator_left_tc__width_512__rotation_1024 (.start(start__rotator_left_tc__width_512__rotation_1024));

rotator_left_tc #(.WIDTH(1024), .ROTATION(0)) rotator_left_tc__width_1024__rotation_0 (.start(start__rotator_left_tc__width_1024__rotation_0));
rotator_left_tc #(.WIDTH(1024), .ROTATION(1)) rotator_left_tc__width_1024__rotation_1 (.start(start__rotator_left_tc__width_1024__rotation_1));
rotator_left_tc #(.WIDTH(1024), .ROTATION(2)) rotator_left_tc__width_1024__rotation_2 (.start(start__rotator_left_tc__width_1024__rotation_2));
rotator_left_tc #(.WIDTH(1024), .ROTATION(3)) rotator_left_tc__width_1024__rotation_3 (.start(start__rotator_left_tc__width_1024__rotation_3));
rotator_left_tc #(.WIDTH(1024), .ROTATION(4)) rotator_left_tc__width_1024__rotation_4 (.start(start__rotator_left_tc__width_1024__rotation_4));
rotator_left_tc #(.WIDTH(1024), .ROTATION(5)) rotator_left_tc__width_1024__rotation_5 (.start(start__rotator_left_tc__width_1024__rotation_5));
rotator_left_tc #(.WIDTH(1024), .ROTATION(6)) rotator_left_tc__width_1024__rotation_6 (.start(start__rotator_left_tc__width_1024__rotation_6));
rotator_left_tc #(.WIDTH(1024), .ROTATION(7)) rotator_left_tc__width_1024__rotation_7 (.start(start__rotator_left_tc__width_1024__rotation_7));
rotator_left_tc #(.WIDTH(1024), .ROTATION(512)) rotator_left_tc__width_1024__rotation_512 (.start(start__rotator_left_tc__width_1024__rotation_512));
rotator_left_tc #(.WIDTH(1024), .ROTATION(1023)) rotator_left_tc__width_1024__rotation_1023 (.start(start__rotator_left_tc__width_1024__rotation_1023));
rotator_left_tc #(.WIDTH(1024), .ROTATION(1024)) rotator_left_tc__width_1024__rotation_1024 (.start(start__rotator_left_tc__width_1024__rotation_1024));
rotator_left_tc #(.WIDTH(1024), .ROTATION(1025)) rotator_left_tc__width_1024__rotation_1025 (.start(start__rotator_left_tc__width_1024__rotation_1025));
rotator_left_tc #(.WIDTH(1024), .ROTATION(1536)) rotator_left_tc__width_1024__rotation_1536 (.start(start__rotator_left_tc__width_1024__rotation_1536));
rotator_left_tc #(.WIDTH(1024), .ROTATION(2047)) rotator_left_tc__width_1024__rotation_2047 (.start(start__rotator_left_tc__width_1024__rotation_2047));
rotator_left_tc #(.WIDTH(1024), .ROTATION(2048)) rotator_left_tc__width_1024__rotation_2048 (.start(start__rotator_left_tc__width_1024__rotation_2048));


initial begin
  // Log waves
  $dumpfile("rotator_left.tb.vcd");
  $dumpvars(0,rotator_left_tc__width_1__rotation_0);
  $dumpvars(0,rotator_left_tc__width_1__rotation_1);

  $dumpvars(0,rotator_left_tc__width_2__rotation_0);
  $dumpvars(0,rotator_left_tc__width_2__rotation_1);
  $dumpvars(0,rotator_left_tc__width_2__rotation_2);
  $dumpvars(0,rotator_left_tc__width_2__rotation_3);

  $dumpvars(0,rotator_left_tc__width_3__rotation_0);
  $dumpvars(0,rotator_left_tc__width_3__rotation_1);
  $dumpvars(0,rotator_left_tc__width_3__rotation_2);
  $dumpvars(0,rotator_left_tc__width_3__rotation_3);
  $dumpvars(0,rotator_left_tc__width_3__rotation_4);
  $dumpvars(0,rotator_left_tc__width_3__rotation_5);

  $dumpvars(0,rotator_left_tc__width_4__rotation_0);
  $dumpvars(0,rotator_left_tc__width_4__rotation_1);
  $dumpvars(0,rotator_left_tc__width_4__rotation_2);
  $dumpvars(0,rotator_left_tc__width_4__rotation_3);
  $dumpvars(0,rotator_left_tc__width_4__rotation_4);
  $dumpvars(0,rotator_left_tc__width_4__rotation_5);
  $dumpvars(0,rotator_left_tc__width_4__rotation_6);
  $dumpvars(0,rotator_left_tc__width_4__rotation_7);

  $dumpvars(0,rotator_left_tc__width_5__rotation_0);
  $dumpvars(0,rotator_left_tc__width_5__rotation_1);
  $dumpvars(0,rotator_left_tc__width_5__rotation_2);
  $dumpvars(0,rotator_left_tc__width_5__rotation_3);
  $dumpvars(0,rotator_left_tc__width_5__rotation_4);
  $dumpvars(0,rotator_left_tc__width_5__rotation_5);
  $dumpvars(0,rotator_left_tc__width_5__rotation_6);
  $dumpvars(0,rotator_left_tc__width_5__rotation_7);
  $dumpvars(0,rotator_left_tc__width_5__rotation_8);
  $dumpvars(0,rotator_left_tc__width_5__rotation_9);

  $dumpvars(0,rotator_left_tc__width_6__rotation_0);
  $dumpvars(0,rotator_left_tc__width_6__rotation_1);
  $dumpvars(0,rotator_left_tc__width_6__rotation_2);
  $dumpvars(0,rotator_left_tc__width_6__rotation_3);
  $dumpvars(0,rotator_left_tc__width_6__rotation_4);
  $dumpvars(0,rotator_left_tc__width_6__rotation_5);
  $dumpvars(0,rotator_left_tc__width_6__rotation_6);
  $dumpvars(0,rotator_left_tc__width_6__rotation_7);
  $dumpvars(0,rotator_left_tc__width_6__rotation_8);
  $dumpvars(0,rotator_left_tc__width_6__rotation_9);
  $dumpvars(0,rotator_left_tc__width_6__rotation_10);
  $dumpvars(0,rotator_left_tc__width_6__rotation_11);

  $dumpvars(0,rotator_left_tc__width_7__rotation_0);
  $dumpvars(0,rotator_left_tc__width_7__rotation_1);
  $dumpvars(0,rotator_left_tc__width_7__rotation_2);
  $dumpvars(0,rotator_left_tc__width_7__rotation_3);
  $dumpvars(0,rotator_left_tc__width_7__rotation_4);
  $dumpvars(0,rotator_left_tc__width_7__rotation_5);
  $dumpvars(0,rotator_left_tc__width_7__rotation_6);
  $dumpvars(0,rotator_left_tc__width_7__rotation_7);
  $dumpvars(0,rotator_left_tc__width_7__rotation_8);
  $dumpvars(0,rotator_left_tc__width_7__rotation_9);
  $dumpvars(0,rotator_left_tc__width_7__rotation_10);
  $dumpvars(0,rotator_left_tc__width_7__rotation_11);
  $dumpvars(0,rotator_left_tc__width_7__rotation_12);
  $dumpvars(0,rotator_left_tc__width_7__rotation_13);

  $dumpvars(0,rotator_left_tc__width_8__rotation_0);
  $dumpvars(0,rotator_left_tc__width_8__rotation_1);
  $dumpvars(0,rotator_left_tc__width_8__rotation_2);
  $dumpvars(0,rotator_left_tc__width_8__rotation_3);
  $dumpvars(0,rotator_left_tc__width_8__rotation_4);
  $dumpvars(0,rotator_left_tc__width_8__rotation_5);
  $dumpvars(0,rotator_left_tc__width_8__rotation_6);
  $dumpvars(0,rotator_left_tc__width_8__rotation_7);
  $dumpvars(0,rotator_left_tc__width_8__rotation_8);
  $dumpvars(0,rotator_left_tc__width_8__rotation_9);
  $dumpvars(0,rotator_left_tc__width_8__rotation_10);
  $dumpvars(0,rotator_left_tc__width_8__rotation_11);
  $dumpvars(0,rotator_left_tc__width_8__rotation_12);
  $dumpvars(0,rotator_left_tc__width_8__rotation_13);
  $dumpvars(0,rotator_left_tc__width_8__rotation_14);
  $dumpvars(0,rotator_left_tc__width_8__rotation_15);

  $dumpvars(0,rotator_left_tc__width_9__rotation_0);
  $dumpvars(0,rotator_left_tc__width_9__rotation_1);
  $dumpvars(0,rotator_left_tc__width_9__rotation_2);
  $dumpvars(0,rotator_left_tc__width_9__rotation_3);
  $dumpvars(0,rotator_left_tc__width_9__rotation_4);
  $dumpvars(0,rotator_left_tc__width_9__rotation_5);
  $dumpvars(0,rotator_left_tc__width_9__rotation_6);
  $dumpvars(0,rotator_left_tc__width_9__rotation_7);
  $dumpvars(0,rotator_left_tc__width_9__rotation_8);
  $dumpvars(0,rotator_left_tc__width_9__rotation_9);
  $dumpvars(0,rotator_left_tc__width_9__rotation_10);
  $dumpvars(0,rotator_left_tc__width_9__rotation_11);
  $dumpvars(0,rotator_left_tc__width_9__rotation_12);
  $dumpvars(0,rotator_left_tc__width_9__rotation_13);
  $dumpvars(0,rotator_left_tc__width_9__rotation_14);
  $dumpvars(0,rotator_left_tc__width_9__rotation_15);
  $dumpvars(0,rotator_left_tc__width_9__rotation_16);
  $dumpvars(0,rotator_left_tc__width_9__rotation_17);

  $dumpvars(0,rotator_left_tc__width_10__rotation_0);
  $dumpvars(0,rotator_left_tc__width_10__rotation_1);
  $dumpvars(0,rotator_left_tc__width_10__rotation_2);
  $dumpvars(0,rotator_left_tc__width_10__rotation_3);
  $dumpvars(0,rotator_left_tc__width_10__rotation_4);
  $dumpvars(0,rotator_left_tc__width_10__rotation_5);
  $dumpvars(0,rotator_left_tc__width_10__rotation_6);
  $dumpvars(0,rotator_left_tc__width_10__rotation_7);
  $dumpvars(0,rotator_left_tc__width_10__rotation_8);
  $dumpvars(0,rotator_left_tc__width_10__rotation_9);
  $dumpvars(0,rotator_left_tc__width_10__rotation_10);
  $dumpvars(0,rotator_left_tc__width_10__rotation_11);
  $dumpvars(0,rotator_left_tc__width_10__rotation_12);
  $dumpvars(0,rotator_left_tc__width_10__rotation_13);
  $dumpvars(0,rotator_left_tc__width_10__rotation_14);
  $dumpvars(0,rotator_left_tc__width_10__rotation_15);
  $dumpvars(0,rotator_left_tc__width_10__rotation_16);
  $dumpvars(0,rotator_left_tc__width_10__rotation_17);
  $dumpvars(0,rotator_left_tc__width_10__rotation_18);
  $dumpvars(0,rotator_left_tc__width_10__rotation_19);

  $dumpvars(0,rotator_left_tc__width_11__rotation_0);
  $dumpvars(0,rotator_left_tc__width_11__rotation_1);
  $dumpvars(0,rotator_left_tc__width_11__rotation_2);
  $dumpvars(0,rotator_left_tc__width_11__rotation_3);
  $dumpvars(0,rotator_left_tc__width_11__rotation_4);
  $dumpvars(0,rotator_left_tc__width_11__rotation_5);
  $dumpvars(0,rotator_left_tc__width_11__rotation_6);
  $dumpvars(0,rotator_left_tc__width_11__rotation_7);
  $dumpvars(0,rotator_left_tc__width_11__rotation_8);
  $dumpvars(0,rotator_left_tc__width_11__rotation_9);
  $dumpvars(0,rotator_left_tc__width_11__rotation_10);
  $dumpvars(0,rotator_left_tc__width_11__rotation_11);
  $dumpvars(0,rotator_left_tc__width_11__rotation_12);
  $dumpvars(0,rotator_left_tc__width_11__rotation_13);
  $dumpvars(0,rotator_left_tc__width_11__rotation_14);
  $dumpvars(0,rotator_left_tc__width_11__rotation_15);
  $dumpvars(0,rotator_left_tc__width_11__rotation_16);
  $dumpvars(0,rotator_left_tc__width_11__rotation_17);
  $dumpvars(0,rotator_left_tc__width_11__rotation_18);
  $dumpvars(0,rotator_left_tc__width_11__rotation_19);
  $dumpvars(0,rotator_left_tc__width_11__rotation_20);
  $dumpvars(0,rotator_left_tc__width_11__rotation_21);

  $dumpvars(0,rotator_left_tc__width_12__rotation_0);
  $dumpvars(0,rotator_left_tc__width_12__rotation_1);
  $dumpvars(0,rotator_left_tc__width_12__rotation_2);
  $dumpvars(0,rotator_left_tc__width_12__rotation_3);
  $dumpvars(0,rotator_left_tc__width_12__rotation_4);
  $dumpvars(0,rotator_left_tc__width_12__rotation_5);
  $dumpvars(0,rotator_left_tc__width_12__rotation_6);
  $dumpvars(0,rotator_left_tc__width_12__rotation_7);
  $dumpvars(0,rotator_left_tc__width_12__rotation_8);
  $dumpvars(0,rotator_left_tc__width_12__rotation_9);
  $dumpvars(0,rotator_left_tc__width_12__rotation_10);
  $dumpvars(0,rotator_left_tc__width_12__rotation_11);
  $dumpvars(0,rotator_left_tc__width_12__rotation_12);
  $dumpvars(0,rotator_left_tc__width_12__rotation_13);
  $dumpvars(0,rotator_left_tc__width_12__rotation_14);
  $dumpvars(0,rotator_left_tc__width_12__rotation_15);
  $dumpvars(0,rotator_left_tc__width_12__rotation_16);
  $dumpvars(0,rotator_left_tc__width_12__rotation_17);
  $dumpvars(0,rotator_left_tc__width_12__rotation_18);
  $dumpvars(0,rotator_left_tc__width_12__rotation_19);
  $dumpvars(0,rotator_left_tc__width_12__rotation_20);
  $dumpvars(0,rotator_left_tc__width_12__rotation_21);
  $dumpvars(0,rotator_left_tc__width_12__rotation_22);
  $dumpvars(0,rotator_left_tc__width_12__rotation_23);

  $dumpvars(0,rotator_left_tc__width_16__rotation_0);
  $dumpvars(0,rotator_left_tc__width_16__rotation_1);
  $dumpvars(0,rotator_left_tc__width_16__rotation_2);
  $dumpvars(0,rotator_left_tc__width_16__rotation_3);
  $dumpvars(0,rotator_left_tc__width_16__rotation_4);
  $dumpvars(0,rotator_left_tc__width_16__rotation_5);
  $dumpvars(0,rotator_left_tc__width_16__rotation_6);
  $dumpvars(0,rotator_left_tc__width_16__rotation_7);
  $dumpvars(0,rotator_left_tc__width_16__rotation_8);
  $dumpvars(0,rotator_left_tc__width_16__rotation_15);
  $dumpvars(0,rotator_left_tc__width_16__rotation_16);
  $dumpvars(0,rotator_left_tc__width_16__rotation_17);
  $dumpvars(0,rotator_left_tc__width_16__rotation_24);
  $dumpvars(0,rotator_left_tc__width_16__rotation_31);
  $dumpvars(0,rotator_left_tc__width_16__rotation_32);

  $dumpvars(0,rotator_left_tc__width_24__rotation_0);
  $dumpvars(0,rotator_left_tc__width_24__rotation_1);
  $dumpvars(0,rotator_left_tc__width_24__rotation_2);
  $dumpvars(0,rotator_left_tc__width_24__rotation_3);
  $dumpvars(0,rotator_left_tc__width_24__rotation_4);
  $dumpvars(0,rotator_left_tc__width_24__rotation_5);
  $dumpvars(0,rotator_left_tc__width_24__rotation_6);
  $dumpvars(0,rotator_left_tc__width_24__rotation_7);
  $dumpvars(0,rotator_left_tc__width_24__rotation_12);
  $dumpvars(0,rotator_left_tc__width_24__rotation_23);
  $dumpvars(0,rotator_left_tc__width_24__rotation_24);
  $dumpvars(0,rotator_left_tc__width_24__rotation_25);
  $dumpvars(0,rotator_left_tc__width_24__rotation_36);
  $dumpvars(0,rotator_left_tc__width_24__rotation_47);
  $dumpvars(0,rotator_left_tc__width_24__rotation_48);

  $dumpvars(0,rotator_left_tc__width_32__rotation_0);
  $dumpvars(0,rotator_left_tc__width_32__rotation_1);
  $dumpvars(0,rotator_left_tc__width_32__rotation_2);
  $dumpvars(0,rotator_left_tc__width_32__rotation_3);
  $dumpvars(0,rotator_left_tc__width_32__rotation_4);
  $dumpvars(0,rotator_left_tc__width_32__rotation_5);
  $dumpvars(0,rotator_left_tc__width_32__rotation_6);
  $dumpvars(0,rotator_left_tc__width_32__rotation_7);
  $dumpvars(0,rotator_left_tc__width_32__rotation_16);
  $dumpvars(0,rotator_left_tc__width_32__rotation_31);
  $dumpvars(0,rotator_left_tc__width_32__rotation_32);
  $dumpvars(0,rotator_left_tc__width_32__rotation_33);
  $dumpvars(0,rotator_left_tc__width_32__rotation_48);
  $dumpvars(0,rotator_left_tc__width_32__rotation_63);
  $dumpvars(0,rotator_left_tc__width_32__rotation_64);

  $dumpvars(0,rotator_left_tc__width_48__rotation_0);
  $dumpvars(0,rotator_left_tc__width_48__rotation_1);
  $dumpvars(0,rotator_left_tc__width_48__rotation_2);
  $dumpvars(0,rotator_left_tc__width_48__rotation_3);
  $dumpvars(0,rotator_left_tc__width_48__rotation_4);
  $dumpvars(0,rotator_left_tc__width_48__rotation_5);
  $dumpvars(0,rotator_left_tc__width_48__rotation_6);
  $dumpvars(0,rotator_left_tc__width_48__rotation_7);
  $dumpvars(0,rotator_left_tc__width_48__rotation_24);
  $dumpvars(0,rotator_left_tc__width_48__rotation_47);
  $dumpvars(0,rotator_left_tc__width_48__rotation_48);
  $dumpvars(0,rotator_left_tc__width_48__rotation_49);
  $dumpvars(0,rotator_left_tc__width_48__rotation_72);
  $dumpvars(0,rotator_left_tc__width_48__rotation_95);
  $dumpvars(0,rotator_left_tc__width_48__rotation_96);

  $dumpvars(0,rotator_left_tc__width_64__rotation_0);
  $dumpvars(0,rotator_left_tc__width_64__rotation_1);
  $dumpvars(0,rotator_left_tc__width_64__rotation_2);
  $dumpvars(0,rotator_left_tc__width_64__rotation_3);
  $dumpvars(0,rotator_left_tc__width_64__rotation_4);
  $dumpvars(0,rotator_left_tc__width_64__rotation_5);
  $dumpvars(0,rotator_left_tc__width_64__rotation_6);
  $dumpvars(0,rotator_left_tc__width_64__rotation_7);
  $dumpvars(0,rotator_left_tc__width_64__rotation_32);
  $dumpvars(0,rotator_left_tc__width_64__rotation_63);
  $dumpvars(0,rotator_left_tc__width_64__rotation_64);
  $dumpvars(0,rotator_left_tc__width_64__rotation_65);
  $dumpvars(0,rotator_left_tc__width_64__rotation_96);
  $dumpvars(0,rotator_left_tc__width_64__rotation_127);
  $dumpvars(0,rotator_left_tc__width_64__rotation_128);

  $dumpvars(0,rotator_left_tc__width_128__rotation_0);
  $dumpvars(0,rotator_left_tc__width_128__rotation_1);
  $dumpvars(0,rotator_left_tc__width_128__rotation_2);
  $dumpvars(0,rotator_left_tc__width_128__rotation_3);
  $dumpvars(0,rotator_left_tc__width_128__rotation_4);
  $dumpvars(0,rotator_left_tc__width_128__rotation_5);
  $dumpvars(0,rotator_left_tc__width_128__rotation_6);
  $dumpvars(0,rotator_left_tc__width_128__rotation_7);
  $dumpvars(0,rotator_left_tc__width_128__rotation_64);
  $dumpvars(0,rotator_left_tc__width_128__rotation_127);
  $dumpvars(0,rotator_left_tc__width_128__rotation_128);
  $dumpvars(0,rotator_left_tc__width_128__rotation_129);
  $dumpvars(0,rotator_left_tc__width_128__rotation_192);
  $dumpvars(0,rotator_left_tc__width_128__rotation_255);
  $dumpvars(0,rotator_left_tc__width_128__rotation_256);

  $dumpvars(0,rotator_left_tc__width_256__rotation_0);
  $dumpvars(0,rotator_left_tc__width_256__rotation_1);
  $dumpvars(0,rotator_left_tc__width_256__rotation_2);
  $dumpvars(0,rotator_left_tc__width_256__rotation_3);
  $dumpvars(0,rotator_left_tc__width_256__rotation_4);
  $dumpvars(0,rotator_left_tc__width_256__rotation_5);
  $dumpvars(0,rotator_left_tc__width_256__rotation_6);
  $dumpvars(0,rotator_left_tc__width_256__rotation_7);
  $dumpvars(0,rotator_left_tc__width_256__rotation_128);
  $dumpvars(0,rotator_left_tc__width_256__rotation_255);
  $dumpvars(0,rotator_left_tc__width_256__rotation_256);
  $dumpvars(0,rotator_left_tc__width_256__rotation_257);
  $dumpvars(0,rotator_left_tc__width_256__rotation_384);
  $dumpvars(0,rotator_left_tc__width_256__rotation_511);
  $dumpvars(0,rotator_left_tc__width_256__rotation_512);

  $dumpvars(0,rotator_left_tc__width_512__rotation_0);
  $dumpvars(0,rotator_left_tc__width_512__rotation_1);
  $dumpvars(0,rotator_left_tc__width_512__rotation_2);
  $dumpvars(0,rotator_left_tc__width_512__rotation_3);
  $dumpvars(0,rotator_left_tc__width_512__rotation_4);
  $dumpvars(0,rotator_left_tc__width_512__rotation_5);
  $dumpvars(0,rotator_left_tc__width_512__rotation_6);
  $dumpvars(0,rotator_left_tc__width_512__rotation_7);
  $dumpvars(0,rotator_left_tc__width_512__rotation_256);
  $dumpvars(0,rotator_left_tc__width_512__rotation_511);
  $dumpvars(0,rotator_left_tc__width_512__rotation_512);
  $dumpvars(0,rotator_left_tc__width_512__rotation_513);
  $dumpvars(0,rotator_left_tc__width_512__rotation_768);
  $dumpvars(0,rotator_left_tc__width_512__rotation_1023);
  $dumpvars(0,rotator_left_tc__width_512__rotation_1024);

  $dumpvars(0,rotator_left_tc__width_1024__rotation_0);
  $dumpvars(0,rotator_left_tc__width_1024__rotation_1);
  $dumpvars(0,rotator_left_tc__width_1024__rotation_2);
  $dumpvars(0,rotator_left_tc__width_1024__rotation_3);
  $dumpvars(0,rotator_left_tc__width_1024__rotation_4);
  $dumpvars(0,rotator_left_tc__width_1024__rotation_5);
  $dumpvars(0,rotator_left_tc__width_1024__rotation_6);
  $dumpvars(0,rotator_left_tc__width_1024__rotation_7);
  $dumpvars(0,rotator_left_tc__width_1024__rotation_512);
  $dumpvars(0,rotator_left_tc__width_1024__rotation_1023);
  $dumpvars(0,rotator_left_tc__width_1024__rotation_1024);
  $dumpvars(0,rotator_left_tc__width_1024__rotation_1025);
  $dumpvars(0,rotator_left_tc__width_1024__rotation_1536);
  $dumpvars(0,rotator_left_tc__width_1024__rotation_2047);
  $dumpvars(0,rotator_left_tc__width_1024__rotation_2048);


  // Initialization
  start__rotator_left_tc__width_1__rotation_0 = 0;
  start__rotator_left_tc__width_1__rotation_1 = 0;

  start__rotator_left_tc__width_2__rotation_0 = 0;
  start__rotator_left_tc__width_2__rotation_1 = 0;
  start__rotator_left_tc__width_2__rotation_2 = 0;
  start__rotator_left_tc__width_2__rotation_3 = 0;

  start__rotator_left_tc__width_3__rotation_0 = 0;
  start__rotator_left_tc__width_3__rotation_1 = 0;
  start__rotator_left_tc__width_3__rotation_2 = 0;
  start__rotator_left_tc__width_3__rotation_3 = 0;
  start__rotator_left_tc__width_3__rotation_4 = 0;
  start__rotator_left_tc__width_3__rotation_5 = 0;

  start__rotator_left_tc__width_4__rotation_0 = 0;
  start__rotator_left_tc__width_4__rotation_1 = 0;
  start__rotator_left_tc__width_4__rotation_2 = 0;
  start__rotator_left_tc__width_4__rotation_3 = 0;
  start__rotator_left_tc__width_4__rotation_4 = 0;
  start__rotator_left_tc__width_4__rotation_5 = 0;
  start__rotator_left_tc__width_4__rotation_6 = 0;
  start__rotator_left_tc__width_4__rotation_7 = 0;

  start__rotator_left_tc__width_5__rotation_0 = 0;
  start__rotator_left_tc__width_5__rotation_1 = 0;
  start__rotator_left_tc__width_5__rotation_2 = 0;
  start__rotator_left_tc__width_5__rotation_3 = 0;
  start__rotator_left_tc__width_5__rotation_4 = 0;
  start__rotator_left_tc__width_5__rotation_5 = 0;
  start__rotator_left_tc__width_5__rotation_6 = 0;
  start__rotator_left_tc__width_5__rotation_7 = 0;
  start__rotator_left_tc__width_5__rotation_8 = 0;
  start__rotator_left_tc__width_5__rotation_9 = 0;

  start__rotator_left_tc__width_6__rotation_0 = 0;
  start__rotator_left_tc__width_6__rotation_1 = 0;
  start__rotator_left_tc__width_6__rotation_2 = 0;
  start__rotator_left_tc__width_6__rotation_3 = 0;
  start__rotator_left_tc__width_6__rotation_4 = 0;
  start__rotator_left_tc__width_6__rotation_5 = 0;
  start__rotator_left_tc__width_6__rotation_6 = 0;
  start__rotator_left_tc__width_6__rotation_7 = 0;
  start__rotator_left_tc__width_6__rotation_8 = 0;
  start__rotator_left_tc__width_6__rotation_9 = 0;
  start__rotator_left_tc__width_6__rotation_10 = 0;
  start__rotator_left_tc__width_6__rotation_11 = 0;

  start__rotator_left_tc__width_7__rotation_0 = 0;
  start__rotator_left_tc__width_7__rotation_1 = 0;
  start__rotator_left_tc__width_7__rotation_2 = 0;
  start__rotator_left_tc__width_7__rotation_3 = 0;
  start__rotator_left_tc__width_7__rotation_4 = 0;
  start__rotator_left_tc__width_7__rotation_5 = 0;
  start__rotator_left_tc__width_7__rotation_6 = 0;
  start__rotator_left_tc__width_7__rotation_7 = 0;
  start__rotator_left_tc__width_7__rotation_8 = 0;
  start__rotator_left_tc__width_7__rotation_9 = 0;
  start__rotator_left_tc__width_7__rotation_10 = 0;
  start__rotator_left_tc__width_7__rotation_11 = 0;
  start__rotator_left_tc__width_7__rotation_12 = 0;
  start__rotator_left_tc__width_7__rotation_13 = 0;

  start__rotator_left_tc__width_8__rotation_0 = 0;
  start__rotator_left_tc__width_8__rotation_1 = 0;
  start__rotator_left_tc__width_8__rotation_2 = 0;
  start__rotator_left_tc__width_8__rotation_3 = 0;
  start__rotator_left_tc__width_8__rotation_4 = 0;
  start__rotator_left_tc__width_8__rotation_5 = 0;
  start__rotator_left_tc__width_8__rotation_6 = 0;
  start__rotator_left_tc__width_8__rotation_7 = 0;
  start__rotator_left_tc__width_8__rotation_8 = 0;
  start__rotator_left_tc__width_8__rotation_9 = 0;
  start__rotator_left_tc__width_8__rotation_10 = 0;
  start__rotator_left_tc__width_8__rotation_11 = 0;
  start__rotator_left_tc__width_8__rotation_12 = 0;
  start__rotator_left_tc__width_8__rotation_13 = 0;
  start__rotator_left_tc__width_8__rotation_14 = 0;
  start__rotator_left_tc__width_8__rotation_15 = 0;

  start__rotator_left_tc__width_9__rotation_0 = 0;
  start__rotator_left_tc__width_9__rotation_1 = 0;
  start__rotator_left_tc__width_9__rotation_2 = 0;
  start__rotator_left_tc__width_9__rotation_3 = 0;
  start__rotator_left_tc__width_9__rotation_4 = 0;
  start__rotator_left_tc__width_9__rotation_5 = 0;
  start__rotator_left_tc__width_9__rotation_6 = 0;
  start__rotator_left_tc__width_9__rotation_7 = 0;
  start__rotator_left_tc__width_9__rotation_8 = 0;
  start__rotator_left_tc__width_9__rotation_9 = 0;
  start__rotator_left_tc__width_9__rotation_10 = 0;
  start__rotator_left_tc__width_9__rotation_11 = 0;
  start__rotator_left_tc__width_9__rotation_12 = 0;
  start__rotator_left_tc__width_9__rotation_13 = 0;
  start__rotator_left_tc__width_9__rotation_14 = 0;
  start__rotator_left_tc__width_9__rotation_15 = 0;
  start__rotator_left_tc__width_9__rotation_16 = 0;
  start__rotator_left_tc__width_9__rotation_17 = 0;

  start__rotator_left_tc__width_10__rotation_0 = 0;
  start__rotator_left_tc__width_10__rotation_1 = 0;
  start__rotator_left_tc__width_10__rotation_2 = 0;
  start__rotator_left_tc__width_10__rotation_3 = 0;
  start__rotator_left_tc__width_10__rotation_4 = 0;
  start__rotator_left_tc__width_10__rotation_5 = 0;
  start__rotator_left_tc__width_10__rotation_6 = 0;
  start__rotator_left_tc__width_10__rotation_7 = 0;
  start__rotator_left_tc__width_10__rotation_8 = 0;
  start__rotator_left_tc__width_10__rotation_9 = 0;
  start__rotator_left_tc__width_10__rotation_10 = 0;
  start__rotator_left_tc__width_10__rotation_11 = 0;
  start__rotator_left_tc__width_10__rotation_12 = 0;
  start__rotator_left_tc__width_10__rotation_13 = 0;
  start__rotator_left_tc__width_10__rotation_14 = 0;
  start__rotator_left_tc__width_10__rotation_15 = 0;
  start__rotator_left_tc__width_10__rotation_16 = 0;
  start__rotator_left_tc__width_10__rotation_17 = 0;
  start__rotator_left_tc__width_10__rotation_18 = 0;
  start__rotator_left_tc__width_10__rotation_19 = 0;

  start__rotator_left_tc__width_11__rotation_0 = 0;
  start__rotator_left_tc__width_11__rotation_1 = 0;
  start__rotator_left_tc__width_11__rotation_2 = 0;
  start__rotator_left_tc__width_11__rotation_3 = 0;
  start__rotator_left_tc__width_11__rotation_4 = 0;
  start__rotator_left_tc__width_11__rotation_5 = 0;
  start__rotator_left_tc__width_11__rotation_6 = 0;
  start__rotator_left_tc__width_11__rotation_7 = 0;
  start__rotator_left_tc__width_11__rotation_8 = 0;
  start__rotator_left_tc__width_11__rotation_9 = 0;
  start__rotator_left_tc__width_11__rotation_10 = 0;
  start__rotator_left_tc__width_11__rotation_11 = 0;
  start__rotator_left_tc__width_11__rotation_12 = 0;
  start__rotator_left_tc__width_11__rotation_13 = 0;
  start__rotator_left_tc__width_11__rotation_14 = 0;
  start__rotator_left_tc__width_11__rotation_15 = 0;
  start__rotator_left_tc__width_11__rotation_16 = 0;
  start__rotator_left_tc__width_11__rotation_17 = 0;
  start__rotator_left_tc__width_11__rotation_18 = 0;
  start__rotator_left_tc__width_11__rotation_19 = 0;
  start__rotator_left_tc__width_11__rotation_20 = 0;
  start__rotator_left_tc__width_11__rotation_21 = 0;

  start__rotator_left_tc__width_12__rotation_0 = 0;
  start__rotator_left_tc__width_12__rotation_1 = 0;
  start__rotator_left_tc__width_12__rotation_2 = 0;
  start__rotator_left_tc__width_12__rotation_3 = 0;
  start__rotator_left_tc__width_12__rotation_4 = 0;
  start__rotator_left_tc__width_12__rotation_5 = 0;
  start__rotator_left_tc__width_12__rotation_6 = 0;
  start__rotator_left_tc__width_12__rotation_7 = 0;
  start__rotator_left_tc__width_12__rotation_8 = 0;
  start__rotator_left_tc__width_12__rotation_9 = 0;
  start__rotator_left_tc__width_12__rotation_10 = 0;
  start__rotator_left_tc__width_12__rotation_11 = 0;
  start__rotator_left_tc__width_12__rotation_12 = 0;
  start__rotator_left_tc__width_12__rotation_13 = 0;
  start__rotator_left_tc__width_12__rotation_14 = 0;
  start__rotator_left_tc__width_12__rotation_15 = 0;
  start__rotator_left_tc__width_12__rotation_16 = 0;
  start__rotator_left_tc__width_12__rotation_17 = 0;
  start__rotator_left_tc__width_12__rotation_18 = 0;
  start__rotator_left_tc__width_12__rotation_19 = 0;
  start__rotator_left_tc__width_12__rotation_20 = 0;
  start__rotator_left_tc__width_12__rotation_21 = 0;
  start__rotator_left_tc__width_12__rotation_22 = 0;
  start__rotator_left_tc__width_12__rotation_23 = 0;

  start__rotator_left_tc__width_16__rotation_0 = 0;
  start__rotator_left_tc__width_16__rotation_1 = 0;
  start__rotator_left_tc__width_16__rotation_2 = 0;
  start__rotator_left_tc__width_16__rotation_3 = 0;
  start__rotator_left_tc__width_16__rotation_4 = 0;
  start__rotator_left_tc__width_16__rotation_5 = 0;
  start__rotator_left_tc__width_16__rotation_6 = 0;
  start__rotator_left_tc__width_16__rotation_7 = 0;
  start__rotator_left_tc__width_16__rotation_8 = 0;
  start__rotator_left_tc__width_16__rotation_15 = 0;
  start__rotator_left_tc__width_16__rotation_16 = 0;
  start__rotator_left_tc__width_16__rotation_17 = 0;
  start__rotator_left_tc__width_16__rotation_24 = 0;
  start__rotator_left_tc__width_16__rotation_31 = 0;
  start__rotator_left_tc__width_16__rotation_32 = 0;

  start__rotator_left_tc__width_24__rotation_0 = 0;
  start__rotator_left_tc__width_24__rotation_1 = 0;
  start__rotator_left_tc__width_24__rotation_2 = 0;
  start__rotator_left_tc__width_24__rotation_3 = 0;
  start__rotator_left_tc__width_24__rotation_4 = 0;
  start__rotator_left_tc__width_24__rotation_5 = 0;
  start__rotator_left_tc__width_24__rotation_6 = 0;
  start__rotator_left_tc__width_24__rotation_7 = 0;
  start__rotator_left_tc__width_24__rotation_12 = 0;
  start__rotator_left_tc__width_24__rotation_23 = 0;
  start__rotator_left_tc__width_24__rotation_24 = 0;
  start__rotator_left_tc__width_24__rotation_25 = 0;
  start__rotator_left_tc__width_24__rotation_36 = 0;
  start__rotator_left_tc__width_24__rotation_47 = 0;
  start__rotator_left_tc__width_24__rotation_48 = 0;

  start__rotator_left_tc__width_32__rotation_0 = 0;
  start__rotator_left_tc__width_32__rotation_1 = 0;
  start__rotator_left_tc__width_32__rotation_2 = 0;
  start__rotator_left_tc__width_32__rotation_3 = 0;
  start__rotator_left_tc__width_32__rotation_4 = 0;
  start__rotator_left_tc__width_32__rotation_5 = 0;
  start__rotator_left_tc__width_32__rotation_6 = 0;
  start__rotator_left_tc__width_32__rotation_7 = 0;
  start__rotator_left_tc__width_32__rotation_16 = 0;
  start__rotator_left_tc__width_32__rotation_31 = 0;
  start__rotator_left_tc__width_32__rotation_32 = 0;
  start__rotator_left_tc__width_32__rotation_33 = 0;
  start__rotator_left_tc__width_32__rotation_48 = 0;
  start__rotator_left_tc__width_32__rotation_63 = 0;
  start__rotator_left_tc__width_32__rotation_64 = 0;

  start__rotator_left_tc__width_48__rotation_0 = 0;
  start__rotator_left_tc__width_48__rotation_1 = 0;
  start__rotator_left_tc__width_48__rotation_2 = 0;
  start__rotator_left_tc__width_48__rotation_3 = 0;
  start__rotator_left_tc__width_48__rotation_4 = 0;
  start__rotator_left_tc__width_48__rotation_5 = 0;
  start__rotator_left_tc__width_48__rotation_6 = 0;
  start__rotator_left_tc__width_48__rotation_7 = 0;
  start__rotator_left_tc__width_48__rotation_24 = 0;
  start__rotator_left_tc__width_48__rotation_47 = 0;
  start__rotator_left_tc__width_48__rotation_48 = 0;
  start__rotator_left_tc__width_48__rotation_49 = 0;
  start__rotator_left_tc__width_48__rotation_72 = 0;
  start__rotator_left_tc__width_48__rotation_95 = 0;
  start__rotator_left_tc__width_48__rotation_96 = 0;

  start__rotator_left_tc__width_64__rotation_0 = 0;
  start__rotator_left_tc__width_64__rotation_1 = 0;
  start__rotator_left_tc__width_64__rotation_2 = 0;
  start__rotator_left_tc__width_64__rotation_3 = 0;
  start__rotator_left_tc__width_64__rotation_4 = 0;
  start__rotator_left_tc__width_64__rotation_5 = 0;
  start__rotator_left_tc__width_64__rotation_6 = 0;
  start__rotator_left_tc__width_64__rotation_7 = 0;
  start__rotator_left_tc__width_64__rotation_32 = 0;
  start__rotator_left_tc__width_64__rotation_63 = 0;
  start__rotator_left_tc__width_64__rotation_64 = 0;
  start__rotator_left_tc__width_64__rotation_65 = 0;
  start__rotator_left_tc__width_64__rotation_96 = 0;
  start__rotator_left_tc__width_64__rotation_127 = 0;
  start__rotator_left_tc__width_64__rotation_128 = 0;

  start__rotator_left_tc__width_128__rotation_0 = 0;
  start__rotator_left_tc__width_128__rotation_1 = 0;
  start__rotator_left_tc__width_128__rotation_2 = 0;
  start__rotator_left_tc__width_128__rotation_3 = 0;
  start__rotator_left_tc__width_128__rotation_4 = 0;
  start__rotator_left_tc__width_128__rotation_5 = 0;
  start__rotator_left_tc__width_128__rotation_6 = 0;
  start__rotator_left_tc__width_128__rotation_7 = 0;
  start__rotator_left_tc__width_128__rotation_64 = 0;
  start__rotator_left_tc__width_128__rotation_127 = 0;
  start__rotator_left_tc__width_128__rotation_128 = 0;
  start__rotator_left_tc__width_128__rotation_129 = 0;
  start__rotator_left_tc__width_128__rotation_192 = 0;
  start__rotator_left_tc__width_128__rotation_255 = 0;
  start__rotator_left_tc__width_128__rotation_256 = 0;

  start__rotator_left_tc__width_256__rotation_0 = 0;
  start__rotator_left_tc__width_256__rotation_1 = 0;
  start__rotator_left_tc__width_256__rotation_2 = 0;
  start__rotator_left_tc__width_256__rotation_3 = 0;
  start__rotator_left_tc__width_256__rotation_4 = 0;
  start__rotator_left_tc__width_256__rotation_5 = 0;
  start__rotator_left_tc__width_256__rotation_6 = 0;
  start__rotator_left_tc__width_256__rotation_7 = 0;
  start__rotator_left_tc__width_256__rotation_128 = 0;
  start__rotator_left_tc__width_256__rotation_255 = 0;
  start__rotator_left_tc__width_256__rotation_256 = 0;
  start__rotator_left_tc__width_256__rotation_257 = 0;
  start__rotator_left_tc__width_256__rotation_384 = 0;
  start__rotator_left_tc__width_256__rotation_511 = 0;
  start__rotator_left_tc__width_256__rotation_512 = 0;

  start__rotator_left_tc__width_512__rotation_0 = 0;
  start__rotator_left_tc__width_512__rotation_1 = 0;
  start__rotator_left_tc__width_512__rotation_2 = 0;
  start__rotator_left_tc__width_512__rotation_3 = 0;
  start__rotator_left_tc__width_512__rotation_4 = 0;
  start__rotator_left_tc__width_512__rotation_5 = 0;
  start__rotator_left_tc__width_512__rotation_6 = 0;
  start__rotator_left_tc__width_512__rotation_7 = 0;
  start__rotator_left_tc__width_512__rotation_256 = 0;
  start__rotator_left_tc__width_512__rotation_511 = 0;
  start__rotator_left_tc__width_512__rotation_512 = 0;
  start__rotator_left_tc__width_512__rotation_513 = 0;
  start__rotator_left_tc__width_512__rotation_768 = 0;
  start__rotator_left_tc__width_512__rotation_1023 = 0;
  start__rotator_left_tc__width_512__rotation_1024 = 0;

  start__rotator_left_tc__width_1024__rotation_0 = 0;
  start__rotator_left_tc__width_1024__rotation_1 = 0;
  start__rotator_left_tc__width_1024__rotation_2 = 0;
  start__rotator_left_tc__width_1024__rotation_3 = 0;
  start__rotator_left_tc__width_1024__rotation_4 = 0;
  start__rotator_left_tc__width_1024__rotation_5 = 0;
  start__rotator_left_tc__width_1024__rotation_6 = 0;
  start__rotator_left_tc__width_1024__rotation_7 = 0;
  start__rotator_left_tc__width_1024__rotation_512 = 0;
  start__rotator_left_tc__width_1024__rotation_1023 = 0;
  start__rotator_left_tc__width_1024__rotation_1024 = 0;
  start__rotator_left_tc__width_1024__rotation_1025 = 0;
  start__rotator_left_tc__width_1024__rotation_1536 = 0;
  start__rotator_left_tc__width_1024__rotation_2047 = 0;
  start__rotator_left_tc__width_1024__rotation_2048 = 0;


  // Start testbenches
  start__rotator_left_tc__width_1__rotation_0 = 1;
  while(!rotator_left_tc__width_1__rotation_0.finished) #(1);
  start__rotator_left_tc__width_1__rotation_1 = 1;
  while(!rotator_left_tc__width_1__rotation_1.finished) #(1);

  start__rotator_left_tc__width_2__rotation_0 = 1;
  while(!rotator_left_tc__width_2__rotation_0.finished) #(1);
  start__rotator_left_tc__width_2__rotation_1 = 1;
  while(!rotator_left_tc__width_2__rotation_1.finished) #(1);
  start__rotator_left_tc__width_2__rotation_2 = 1;
  while(!rotator_left_tc__width_2__rotation_2.finished) #(1);
  start__rotator_left_tc__width_2__rotation_3 = 1;
  while(!rotator_left_tc__width_2__rotation_3.finished) #(1);

  start__rotator_left_tc__width_3__rotation_0 = 1;
  while(!rotator_left_tc__width_3__rotation_0.finished) #(1);
  start__rotator_left_tc__width_3__rotation_1 = 1;
  while(!rotator_left_tc__width_3__rotation_1.finished) #(1);
  start__rotator_left_tc__width_3__rotation_2 = 1;
  while(!rotator_left_tc__width_3__rotation_2.finished) #(1);
  start__rotator_left_tc__width_3__rotation_3 = 1;
  while(!rotator_left_tc__width_3__rotation_3.finished) #(1);
  start__rotator_left_tc__width_3__rotation_4 = 1;
  while(!rotator_left_tc__width_3__rotation_4.finished) #(1);
  start__rotator_left_tc__width_3__rotation_5 = 1;
  while(!rotator_left_tc__width_3__rotation_5.finished) #(1);

  start__rotator_left_tc__width_4__rotation_0 = 1;
  while(!rotator_left_tc__width_4__rotation_0.finished) #(1);
  start__rotator_left_tc__width_4__rotation_1 = 1;
  while(!rotator_left_tc__width_4__rotation_1.finished) #(1);
  start__rotator_left_tc__width_4__rotation_2 = 1;
  while(!rotator_left_tc__width_4__rotation_2.finished) #(1);
  start__rotator_left_tc__width_4__rotation_3 = 1;
  while(!rotator_left_tc__width_4__rotation_3.finished) #(1);
  start__rotator_left_tc__width_4__rotation_4 = 1;
  while(!rotator_left_tc__width_4__rotation_4.finished) #(1);
  start__rotator_left_tc__width_4__rotation_5 = 1;
  while(!rotator_left_tc__width_4__rotation_5.finished) #(1);
  start__rotator_left_tc__width_4__rotation_6 = 1;
  while(!rotator_left_tc__width_4__rotation_6.finished) #(1);
  start__rotator_left_tc__width_4__rotation_7 = 1;
  while(!rotator_left_tc__width_4__rotation_7.finished) #(1);

  start__rotator_left_tc__width_5__rotation_0 = 1;
  while(!rotator_left_tc__width_5__rotation_0.finished) #(1);
  start__rotator_left_tc__width_5__rotation_1 = 1;
  while(!rotator_left_tc__width_5__rotation_1.finished) #(1);
  start__rotator_left_tc__width_5__rotation_2 = 1;
  while(!rotator_left_tc__width_5__rotation_2.finished) #(1);
  start__rotator_left_tc__width_5__rotation_3 = 1;
  while(!rotator_left_tc__width_5__rotation_3.finished) #(1);
  start__rotator_left_tc__width_5__rotation_4 = 1;
  while(!rotator_left_tc__width_5__rotation_4.finished) #(1);
  start__rotator_left_tc__width_5__rotation_5 = 1;
  while(!rotator_left_tc__width_5__rotation_5.finished) #(1);
  start__rotator_left_tc__width_5__rotation_6 = 1;
  while(!rotator_left_tc__width_5__rotation_6.finished) #(1);
  start__rotator_left_tc__width_5__rotation_7 = 1;
  while(!rotator_left_tc__width_5__rotation_7.finished) #(1);
  start__rotator_left_tc__width_5__rotation_8 = 1;
  while(!rotator_left_tc__width_5__rotation_8.finished) #(1);
  start__rotator_left_tc__width_5__rotation_9 = 1;
  while(!rotator_left_tc__width_5__rotation_9.finished) #(1);

  start__rotator_left_tc__width_6__rotation_0 = 1;
  while(!rotator_left_tc__width_6__rotation_0.finished) #(1);
  start__rotator_left_tc__width_6__rotation_1 = 1;
  while(!rotator_left_tc__width_6__rotation_1.finished) #(1);
  start__rotator_left_tc__width_6__rotation_2 = 1;
  while(!rotator_left_tc__width_6__rotation_2.finished) #(1);
  start__rotator_left_tc__width_6__rotation_3 = 1;
  while(!rotator_left_tc__width_6__rotation_3.finished) #(1);
  start__rotator_left_tc__width_6__rotation_4 = 1;
  while(!rotator_left_tc__width_6__rotation_4.finished) #(1);
  start__rotator_left_tc__width_6__rotation_5 = 1;
  while(!rotator_left_tc__width_6__rotation_5.finished) #(1);
  start__rotator_left_tc__width_6__rotation_6 = 1;
  while(!rotator_left_tc__width_6__rotation_6.finished) #(1);
  start__rotator_left_tc__width_6__rotation_7 = 1;
  while(!rotator_left_tc__width_6__rotation_7.finished) #(1);
  start__rotator_left_tc__width_6__rotation_8 = 1;
  while(!rotator_left_tc__width_6__rotation_8.finished) #(1);
  start__rotator_left_tc__width_6__rotation_9 = 1;
  while(!rotator_left_tc__width_6__rotation_9.finished) #(1);
  start__rotator_left_tc__width_6__rotation_10 = 1;
  while(!rotator_left_tc__width_6__rotation_10.finished) #(1);
  start__rotator_left_tc__width_6__rotation_11 = 1;
  while(!rotator_left_tc__width_6__rotation_11.finished) #(1);

  start__rotator_left_tc__width_7__rotation_0 = 1;
  while(!rotator_left_tc__width_7__rotation_0.finished) #(1);
  start__rotator_left_tc__width_7__rotation_1 = 1;
  while(!rotator_left_tc__width_7__rotation_1.finished) #(1);
  start__rotator_left_tc__width_7__rotation_2 = 1;
  while(!rotator_left_tc__width_7__rotation_2.finished) #(1);
  start__rotator_left_tc__width_7__rotation_3 = 1;
  while(!rotator_left_tc__width_7__rotation_3.finished) #(1);
  start__rotator_left_tc__width_7__rotation_4 = 1;
  while(!rotator_left_tc__width_7__rotation_4.finished) #(1);
  start__rotator_left_tc__width_7__rotation_5 = 1;
  while(!rotator_left_tc__width_7__rotation_5.finished) #(1);
  start__rotator_left_tc__width_7__rotation_6 = 1;
  while(!rotator_left_tc__width_7__rotation_6.finished) #(1);
  start__rotator_left_tc__width_7__rotation_7 = 1;
  while(!rotator_left_tc__width_7__rotation_7.finished) #(1);
  start__rotator_left_tc__width_7__rotation_8 = 1;
  while(!rotator_left_tc__width_7__rotation_8.finished) #(1);
  start__rotator_left_tc__width_7__rotation_9 = 1;
  while(!rotator_left_tc__width_7__rotation_9.finished) #(1);
  start__rotator_left_tc__width_7__rotation_10 = 1;
  while(!rotator_left_tc__width_7__rotation_10.finished) #(1);
  start__rotator_left_tc__width_7__rotation_11 = 1;
  while(!rotator_left_tc__width_7__rotation_11.finished) #(1);
  start__rotator_left_tc__width_7__rotation_12 = 1;
  while(!rotator_left_tc__width_7__rotation_12.finished) #(1);
  start__rotator_left_tc__width_7__rotation_13 = 1;
  while(!rotator_left_tc__width_7__rotation_13.finished) #(1);

  start__rotator_left_tc__width_8__rotation_0 = 1;
  while(!rotator_left_tc__width_8__rotation_0.finished) #(1);
  start__rotator_left_tc__width_8__rotation_1 = 1;
  while(!rotator_left_tc__width_8__rotation_1.finished) #(1);
  start__rotator_left_tc__width_8__rotation_2 = 1;
  while(!rotator_left_tc__width_8__rotation_2.finished) #(1);
  start__rotator_left_tc__width_8__rotation_3 = 1;
  while(!rotator_left_tc__width_8__rotation_3.finished) #(1);
  start__rotator_left_tc__width_8__rotation_4 = 1;
  while(!rotator_left_tc__width_8__rotation_4.finished) #(1);
  start__rotator_left_tc__width_8__rotation_5 = 1;
  while(!rotator_left_tc__width_8__rotation_5.finished) #(1);
  start__rotator_left_tc__width_8__rotation_6 = 1;
  while(!rotator_left_tc__width_8__rotation_6.finished) #(1);
  start__rotator_left_tc__width_8__rotation_7 = 1;
  while(!rotator_left_tc__width_8__rotation_7.finished) #(1);
  start__rotator_left_tc__width_8__rotation_8 = 1;
  while(!rotator_left_tc__width_8__rotation_8.finished) #(1);
  start__rotator_left_tc__width_8__rotation_9 = 1;
  while(!rotator_left_tc__width_8__rotation_9.finished) #(1);
  start__rotator_left_tc__width_8__rotation_10 = 1;
  while(!rotator_left_tc__width_8__rotation_10.finished) #(1);
  start__rotator_left_tc__width_8__rotation_11 = 1;
  while(!rotator_left_tc__width_8__rotation_11.finished) #(1);
  start__rotator_left_tc__width_8__rotation_12 = 1;
  while(!rotator_left_tc__width_8__rotation_12.finished) #(1);
  start__rotator_left_tc__width_8__rotation_13 = 1;
  while(!rotator_left_tc__width_8__rotation_13.finished) #(1);
  start__rotator_left_tc__width_8__rotation_14 = 1;
  while(!rotator_left_tc__width_8__rotation_14.finished) #(1);
  start__rotator_left_tc__width_8__rotation_15 = 1;
  while(!rotator_left_tc__width_8__rotation_15.finished) #(1);

  start__rotator_left_tc__width_9__rotation_0 = 1;
  while(!rotator_left_tc__width_9__rotation_0.finished) #(1);
  start__rotator_left_tc__width_9__rotation_1 = 1;
  while(!rotator_left_tc__width_9__rotation_1.finished) #(1);
  start__rotator_left_tc__width_9__rotation_2 = 1;
  while(!rotator_left_tc__width_9__rotation_2.finished) #(1);
  start__rotator_left_tc__width_9__rotation_3 = 1;
  while(!rotator_left_tc__width_9__rotation_3.finished) #(1);
  start__rotator_left_tc__width_9__rotation_4 = 1;
  while(!rotator_left_tc__width_9__rotation_4.finished) #(1);
  start__rotator_left_tc__width_9__rotation_5 = 1;
  while(!rotator_left_tc__width_9__rotation_5.finished) #(1);
  start__rotator_left_tc__width_9__rotation_6 = 1;
  while(!rotator_left_tc__width_9__rotation_6.finished) #(1);
  start__rotator_left_tc__width_9__rotation_7 = 1;
  while(!rotator_left_tc__width_9__rotation_7.finished) #(1);
  start__rotator_left_tc__width_9__rotation_8 = 1;
  while(!rotator_left_tc__width_9__rotation_8.finished) #(1);
  start__rotator_left_tc__width_9__rotation_9 = 1;
  while(!rotator_left_tc__width_9__rotation_9.finished) #(1);
  start__rotator_left_tc__width_9__rotation_10 = 1;
  while(!rotator_left_tc__width_9__rotation_10.finished) #(1);
  start__rotator_left_tc__width_9__rotation_11 = 1;
  while(!rotator_left_tc__width_9__rotation_11.finished) #(1);
  start__rotator_left_tc__width_9__rotation_12 = 1;
  while(!rotator_left_tc__width_9__rotation_12.finished) #(1);
  start__rotator_left_tc__width_9__rotation_13 = 1;
  while(!rotator_left_tc__width_9__rotation_13.finished) #(1);
  start__rotator_left_tc__width_9__rotation_14 = 1;
  while(!rotator_left_tc__width_9__rotation_14.finished) #(1);
  start__rotator_left_tc__width_9__rotation_15 = 1;
  while(!rotator_left_tc__width_9__rotation_15.finished) #(1);
  start__rotator_left_tc__width_9__rotation_16 = 1;
  while(!rotator_left_tc__width_9__rotation_16.finished) #(1);
  start__rotator_left_tc__width_9__rotation_17 = 1;
  while(!rotator_left_tc__width_9__rotation_17.finished) #(1);

  start__rotator_left_tc__width_10__rotation_0 = 1;
  while(!rotator_left_tc__width_10__rotation_0.finished) #(1);
  start__rotator_left_tc__width_10__rotation_1 = 1;
  while(!rotator_left_tc__width_10__rotation_1.finished) #(1);
  start__rotator_left_tc__width_10__rotation_2 = 1;
  while(!rotator_left_tc__width_10__rotation_2.finished) #(1);
  start__rotator_left_tc__width_10__rotation_3 = 1;
  while(!rotator_left_tc__width_10__rotation_3.finished) #(1);
  start__rotator_left_tc__width_10__rotation_4 = 1;
  while(!rotator_left_tc__width_10__rotation_4.finished) #(1);
  start__rotator_left_tc__width_10__rotation_5 = 1;
  while(!rotator_left_tc__width_10__rotation_5.finished) #(1);
  start__rotator_left_tc__width_10__rotation_6 = 1;
  while(!rotator_left_tc__width_10__rotation_6.finished) #(1);
  start__rotator_left_tc__width_10__rotation_7 = 1;
  while(!rotator_left_tc__width_10__rotation_7.finished) #(1);
  start__rotator_left_tc__width_10__rotation_8 = 1;
  while(!rotator_left_tc__width_10__rotation_8.finished) #(1);
  start__rotator_left_tc__width_10__rotation_9 = 1;
  while(!rotator_left_tc__width_10__rotation_9.finished) #(1);
  start__rotator_left_tc__width_10__rotation_10 = 1;
  while(!rotator_left_tc__width_10__rotation_10.finished) #(1);
  start__rotator_left_tc__width_10__rotation_11 = 1;
  while(!rotator_left_tc__width_10__rotation_11.finished) #(1);
  start__rotator_left_tc__width_10__rotation_12 = 1;
  while(!rotator_left_tc__width_10__rotation_12.finished) #(1);
  start__rotator_left_tc__width_10__rotation_13 = 1;
  while(!rotator_left_tc__width_10__rotation_13.finished) #(1);
  start__rotator_left_tc__width_10__rotation_14 = 1;
  while(!rotator_left_tc__width_10__rotation_14.finished) #(1);
  start__rotator_left_tc__width_10__rotation_15 = 1;
  while(!rotator_left_tc__width_10__rotation_15.finished) #(1);
  start__rotator_left_tc__width_10__rotation_16 = 1;
  while(!rotator_left_tc__width_10__rotation_16.finished) #(1);
  start__rotator_left_tc__width_10__rotation_17 = 1;
  while(!rotator_left_tc__width_10__rotation_17.finished) #(1);
  start__rotator_left_tc__width_10__rotation_18 = 1;
  while(!rotator_left_tc__width_10__rotation_18.finished) #(1);
  start__rotator_left_tc__width_10__rotation_19 = 1;
  while(!rotator_left_tc__width_10__rotation_19.finished) #(1);

  start__rotator_left_tc__width_11__rotation_0 = 1;
  while(!rotator_left_tc__width_11__rotation_0.finished) #(1);
  start__rotator_left_tc__width_11__rotation_1 = 1;
  while(!rotator_left_tc__width_11__rotation_1.finished) #(1);
  start__rotator_left_tc__width_11__rotation_2 = 1;
  while(!rotator_left_tc__width_11__rotation_2.finished) #(1);
  start__rotator_left_tc__width_11__rotation_3 = 1;
  while(!rotator_left_tc__width_11__rotation_3.finished) #(1);
  start__rotator_left_tc__width_11__rotation_4 = 1;
  while(!rotator_left_tc__width_11__rotation_4.finished) #(1);
  start__rotator_left_tc__width_11__rotation_5 = 1;
  while(!rotator_left_tc__width_11__rotation_5.finished) #(1);
  start__rotator_left_tc__width_11__rotation_6 = 1;
  while(!rotator_left_tc__width_11__rotation_6.finished) #(1);
  start__rotator_left_tc__width_11__rotation_7 = 1;
  while(!rotator_left_tc__width_11__rotation_7.finished) #(1);
  start__rotator_left_tc__width_11__rotation_8 = 1;
  while(!rotator_left_tc__width_11__rotation_8.finished) #(1);
  start__rotator_left_tc__width_11__rotation_9 = 1;
  while(!rotator_left_tc__width_11__rotation_9.finished) #(1);
  start__rotator_left_tc__width_11__rotation_10 = 1;
  while(!rotator_left_tc__width_11__rotation_10.finished) #(1);
  start__rotator_left_tc__width_11__rotation_11 = 1;
  while(!rotator_left_tc__width_11__rotation_11.finished) #(1);
  start__rotator_left_tc__width_11__rotation_12 = 1;
  while(!rotator_left_tc__width_11__rotation_12.finished) #(1);
  start__rotator_left_tc__width_11__rotation_13 = 1;
  while(!rotator_left_tc__width_11__rotation_13.finished) #(1);
  start__rotator_left_tc__width_11__rotation_14 = 1;
  while(!rotator_left_tc__width_11__rotation_14.finished) #(1);
  start__rotator_left_tc__width_11__rotation_15 = 1;
  while(!rotator_left_tc__width_11__rotation_15.finished) #(1);
  start__rotator_left_tc__width_11__rotation_16 = 1;
  while(!rotator_left_tc__width_11__rotation_16.finished) #(1);
  start__rotator_left_tc__width_11__rotation_17 = 1;
  while(!rotator_left_tc__width_11__rotation_17.finished) #(1);
  start__rotator_left_tc__width_11__rotation_18 = 1;
  while(!rotator_left_tc__width_11__rotation_18.finished) #(1);
  start__rotator_left_tc__width_11__rotation_19 = 1;
  while(!rotator_left_tc__width_11__rotation_19.finished) #(1);
  start__rotator_left_tc__width_11__rotation_20 = 1;
  while(!rotator_left_tc__width_11__rotation_20.finished) #(1);
  start__rotator_left_tc__width_11__rotation_21 = 1;
  while(!rotator_left_tc__width_11__rotation_21.finished) #(1);

  start__rotator_left_tc__width_12__rotation_0 = 1;
  while(!rotator_left_tc__width_12__rotation_0.finished) #(1);
  start__rotator_left_tc__width_12__rotation_1 = 1;
  while(!rotator_left_tc__width_12__rotation_1.finished) #(1);
  start__rotator_left_tc__width_12__rotation_2 = 1;
  while(!rotator_left_tc__width_12__rotation_2.finished) #(1);
  start__rotator_left_tc__width_12__rotation_3 = 1;
  while(!rotator_left_tc__width_12__rotation_3.finished) #(1);
  start__rotator_left_tc__width_12__rotation_4 = 1;
  while(!rotator_left_tc__width_12__rotation_4.finished) #(1);
  start__rotator_left_tc__width_12__rotation_5 = 1;
  while(!rotator_left_tc__width_12__rotation_5.finished) #(1);
  start__rotator_left_tc__width_12__rotation_6 = 1;
  while(!rotator_left_tc__width_12__rotation_6.finished) #(1);
  start__rotator_left_tc__width_12__rotation_7 = 1;
  while(!rotator_left_tc__width_12__rotation_7.finished) #(1);
  start__rotator_left_tc__width_12__rotation_8 = 1;
  while(!rotator_left_tc__width_12__rotation_8.finished) #(1);
  start__rotator_left_tc__width_12__rotation_9 = 1;
  while(!rotator_left_tc__width_12__rotation_9.finished) #(1);
  start__rotator_left_tc__width_12__rotation_10 = 1;
  while(!rotator_left_tc__width_12__rotation_10.finished) #(1);
  start__rotator_left_tc__width_12__rotation_11 = 1;
  while(!rotator_left_tc__width_12__rotation_11.finished) #(1);
  start__rotator_left_tc__width_12__rotation_12 = 1;
  while(!rotator_left_tc__width_12__rotation_12.finished) #(1);
  start__rotator_left_tc__width_12__rotation_13 = 1;
  while(!rotator_left_tc__width_12__rotation_13.finished) #(1);
  start__rotator_left_tc__width_12__rotation_14 = 1;
  while(!rotator_left_tc__width_12__rotation_14.finished) #(1);
  start__rotator_left_tc__width_12__rotation_15 = 1;
  while(!rotator_left_tc__width_12__rotation_15.finished) #(1);
  start__rotator_left_tc__width_12__rotation_16 = 1;
  while(!rotator_left_tc__width_12__rotation_16.finished) #(1);
  start__rotator_left_tc__width_12__rotation_17 = 1;
  while(!rotator_left_tc__width_12__rotation_17.finished) #(1);
  start__rotator_left_tc__width_12__rotation_18 = 1;
  while(!rotator_left_tc__width_12__rotation_18.finished) #(1);
  start__rotator_left_tc__width_12__rotation_19 = 1;
  while(!rotator_left_tc__width_12__rotation_19.finished) #(1);
  start__rotator_left_tc__width_12__rotation_20 = 1;
  while(!rotator_left_tc__width_12__rotation_20.finished) #(1);
  start__rotator_left_tc__width_12__rotation_21 = 1;
  while(!rotator_left_tc__width_12__rotation_21.finished) #(1);
  start__rotator_left_tc__width_12__rotation_22 = 1;
  while(!rotator_left_tc__width_12__rotation_22.finished) #(1);
  start__rotator_left_tc__width_12__rotation_23 = 1;
  while(!rotator_left_tc__width_12__rotation_23.finished) #(1);

  start__rotator_left_tc__width_16__rotation_0 = 1;
  while(!rotator_left_tc__width_16__rotation_0.finished) #(1);
  start__rotator_left_tc__width_16__rotation_1 = 1;
  while(!rotator_left_tc__width_16__rotation_1.finished) #(1);
  start__rotator_left_tc__width_16__rotation_2 = 1;
  while(!rotator_left_tc__width_16__rotation_2.finished) #(1);
  start__rotator_left_tc__width_16__rotation_3 = 1;
  while(!rotator_left_tc__width_16__rotation_3.finished) #(1);
  start__rotator_left_tc__width_16__rotation_4 = 1;
  while(!rotator_left_tc__width_16__rotation_4.finished) #(1);
  start__rotator_left_tc__width_16__rotation_5 = 1;
  while(!rotator_left_tc__width_16__rotation_5.finished) #(1);
  start__rotator_left_tc__width_16__rotation_6 = 1;
  while(!rotator_left_tc__width_16__rotation_6.finished) #(1);
  start__rotator_left_tc__width_16__rotation_7 = 1;
  while(!rotator_left_tc__width_16__rotation_7.finished) #(1);
  start__rotator_left_tc__width_16__rotation_8 = 1;
  while(!rotator_left_tc__width_16__rotation_8.finished) #(1);
  start__rotator_left_tc__width_16__rotation_15 = 1;
  while(!rotator_left_tc__width_16__rotation_15.finished) #(1);
  start__rotator_left_tc__width_16__rotation_16 = 1;
  while(!rotator_left_tc__width_16__rotation_16.finished) #(1);
  start__rotator_left_tc__width_16__rotation_17 = 1;
  while(!rotator_left_tc__width_16__rotation_17.finished) #(1);
  start__rotator_left_tc__width_16__rotation_24 = 1;
  while(!rotator_left_tc__width_16__rotation_24.finished) #(1);
  start__rotator_left_tc__width_16__rotation_31 = 1;
  while(!rotator_left_tc__width_16__rotation_31.finished) #(1);
  start__rotator_left_tc__width_16__rotation_32 = 1;
  while(!rotator_left_tc__width_16__rotation_32.finished) #(1);

  start__rotator_left_tc__width_24__rotation_0 = 1;
  while(!rotator_left_tc__width_24__rotation_0.finished) #(1);
  start__rotator_left_tc__width_24__rotation_1 = 1;
  while(!rotator_left_tc__width_24__rotation_1.finished) #(1);
  start__rotator_left_tc__width_24__rotation_2 = 1;
  while(!rotator_left_tc__width_24__rotation_2.finished) #(1);
  start__rotator_left_tc__width_24__rotation_3 = 1;
  while(!rotator_left_tc__width_24__rotation_3.finished) #(1);
  start__rotator_left_tc__width_24__rotation_4 = 1;
  while(!rotator_left_tc__width_24__rotation_4.finished) #(1);
  start__rotator_left_tc__width_24__rotation_5 = 1;
  while(!rotator_left_tc__width_24__rotation_5.finished) #(1);
  start__rotator_left_tc__width_24__rotation_6 = 1;
  while(!rotator_left_tc__width_24__rotation_6.finished) #(1);
  start__rotator_left_tc__width_24__rotation_7 = 1;
  while(!rotator_left_tc__width_24__rotation_7.finished) #(1);
  start__rotator_left_tc__width_24__rotation_12 = 1;
  while(!rotator_left_tc__width_24__rotation_12.finished) #(1);
  start__rotator_left_tc__width_24__rotation_23 = 1;
  while(!rotator_left_tc__width_24__rotation_23.finished) #(1);
  start__rotator_left_tc__width_24__rotation_24 = 1;
  while(!rotator_left_tc__width_24__rotation_24.finished) #(1);
  start__rotator_left_tc__width_24__rotation_25 = 1;
  while(!rotator_left_tc__width_24__rotation_25.finished) #(1);
  start__rotator_left_tc__width_24__rotation_36 = 1;
  while(!rotator_left_tc__width_24__rotation_36.finished) #(1);
  start__rotator_left_tc__width_24__rotation_47 = 1;
  while(!rotator_left_tc__width_24__rotation_47.finished) #(1);
  start__rotator_left_tc__width_24__rotation_48 = 1;
  while(!rotator_left_tc__width_24__rotation_48.finished) #(1);

  start__rotator_left_tc__width_32__rotation_0 = 1;
  while(!rotator_left_tc__width_32__rotation_0.finished) #(1);
  start__rotator_left_tc__width_32__rotation_1 = 1;
  while(!rotator_left_tc__width_32__rotation_1.finished) #(1);
  start__rotator_left_tc__width_32__rotation_2 = 1;
  while(!rotator_left_tc__width_32__rotation_2.finished) #(1);
  start__rotator_left_tc__width_32__rotation_3 = 1;
  while(!rotator_left_tc__width_32__rotation_3.finished) #(1);
  start__rotator_left_tc__width_32__rotation_4 = 1;
  while(!rotator_left_tc__width_32__rotation_4.finished) #(1);
  start__rotator_left_tc__width_32__rotation_5 = 1;
  while(!rotator_left_tc__width_32__rotation_5.finished) #(1);
  start__rotator_left_tc__width_32__rotation_6 = 1;
  while(!rotator_left_tc__width_32__rotation_6.finished) #(1);
  start__rotator_left_tc__width_32__rotation_7 = 1;
  while(!rotator_left_tc__width_32__rotation_7.finished) #(1);
  start__rotator_left_tc__width_32__rotation_16 = 1;
  while(!rotator_left_tc__width_32__rotation_16.finished) #(1);
  start__rotator_left_tc__width_32__rotation_31 = 1;
  while(!rotator_left_tc__width_32__rotation_31.finished) #(1);
  start__rotator_left_tc__width_32__rotation_32 = 1;
  while(!rotator_left_tc__width_32__rotation_32.finished) #(1);
  start__rotator_left_tc__width_32__rotation_33 = 1;
  while(!rotator_left_tc__width_32__rotation_33.finished) #(1);
  start__rotator_left_tc__width_32__rotation_48 = 1;
  while(!rotator_left_tc__width_32__rotation_48.finished) #(1);
  start__rotator_left_tc__width_32__rotation_63 = 1;
  while(!rotator_left_tc__width_32__rotation_63.finished) #(1);
  start__rotator_left_tc__width_32__rotation_64 = 1;
  while(!rotator_left_tc__width_32__rotation_64.finished) #(1);

  start__rotator_left_tc__width_48__rotation_0 = 1;
  while(!rotator_left_tc__width_48__rotation_0.finished) #(1);
  start__rotator_left_tc__width_48__rotation_1 = 1;
  while(!rotator_left_tc__width_48__rotation_1.finished) #(1);
  start__rotator_left_tc__width_48__rotation_2 = 1;
  while(!rotator_left_tc__width_48__rotation_2.finished) #(1);
  start__rotator_left_tc__width_48__rotation_3 = 1;
  while(!rotator_left_tc__width_48__rotation_3.finished) #(1);
  start__rotator_left_tc__width_48__rotation_4 = 1;
  while(!rotator_left_tc__width_48__rotation_4.finished) #(1);
  start__rotator_left_tc__width_48__rotation_5 = 1;
  while(!rotator_left_tc__width_48__rotation_5.finished) #(1);
  start__rotator_left_tc__width_48__rotation_6 = 1;
  while(!rotator_left_tc__width_48__rotation_6.finished) #(1);
  start__rotator_left_tc__width_48__rotation_7 = 1;
  while(!rotator_left_tc__width_48__rotation_7.finished) #(1);
  start__rotator_left_tc__width_48__rotation_24 = 1;
  while(!rotator_left_tc__width_48__rotation_24.finished) #(1);
  start__rotator_left_tc__width_48__rotation_47 = 1;
  while(!rotator_left_tc__width_48__rotation_47.finished) #(1);
  start__rotator_left_tc__width_48__rotation_48 = 1;
  while(!rotator_left_tc__width_48__rotation_48.finished) #(1);
  start__rotator_left_tc__width_48__rotation_49 = 1;
  while(!rotator_left_tc__width_48__rotation_49.finished) #(1);
  start__rotator_left_tc__width_48__rotation_72 = 1;
  while(!rotator_left_tc__width_48__rotation_72.finished) #(1);
  start__rotator_left_tc__width_48__rotation_95 = 1;
  while(!rotator_left_tc__width_48__rotation_95.finished) #(1);
  start__rotator_left_tc__width_48__rotation_96 = 1;
  while(!rotator_left_tc__width_48__rotation_96.finished) #(1);

  start__rotator_left_tc__width_64__rotation_0 = 1;
  while(!rotator_left_tc__width_64__rotation_0.finished) #(1);
  start__rotator_left_tc__width_64__rotation_1 = 1;
  while(!rotator_left_tc__width_64__rotation_1.finished) #(1);
  start__rotator_left_tc__width_64__rotation_2 = 1;
  while(!rotator_left_tc__width_64__rotation_2.finished) #(1);
  start__rotator_left_tc__width_64__rotation_3 = 1;
  while(!rotator_left_tc__width_64__rotation_3.finished) #(1);
  start__rotator_left_tc__width_64__rotation_4 = 1;
  while(!rotator_left_tc__width_64__rotation_4.finished) #(1);
  start__rotator_left_tc__width_64__rotation_5 = 1;
  while(!rotator_left_tc__width_64__rotation_5.finished) #(1);
  start__rotator_left_tc__width_64__rotation_6 = 1;
  while(!rotator_left_tc__width_64__rotation_6.finished) #(1);
  start__rotator_left_tc__width_64__rotation_7 = 1;
  while(!rotator_left_tc__width_64__rotation_7.finished) #(1);
  start__rotator_left_tc__width_64__rotation_32 = 1;
  while(!rotator_left_tc__width_64__rotation_32.finished) #(1);
  start__rotator_left_tc__width_64__rotation_63 = 1;
  while(!rotator_left_tc__width_64__rotation_63.finished) #(1);
  start__rotator_left_tc__width_64__rotation_64 = 1;
  while(!rotator_left_tc__width_64__rotation_64.finished) #(1);
  start__rotator_left_tc__width_64__rotation_65 = 1;
  while(!rotator_left_tc__width_64__rotation_65.finished) #(1);
  start__rotator_left_tc__width_64__rotation_96 = 1;
  while(!rotator_left_tc__width_64__rotation_96.finished) #(1);
  start__rotator_left_tc__width_64__rotation_127 = 1;
  while(!rotator_left_tc__width_64__rotation_127.finished) #(1);
  start__rotator_left_tc__width_64__rotation_128 = 1;
  while(!rotator_left_tc__width_64__rotation_128.finished) #(1);

  start__rotator_left_tc__width_128__rotation_0 = 1;
  while(!rotator_left_tc__width_128__rotation_0.finished) #(1);
  start__rotator_left_tc__width_128__rotation_1 = 1;
  while(!rotator_left_tc__width_128__rotation_1.finished) #(1);
  start__rotator_left_tc__width_128__rotation_2 = 1;
  while(!rotator_left_tc__width_128__rotation_2.finished) #(1);
  start__rotator_left_tc__width_128__rotation_3 = 1;
  while(!rotator_left_tc__width_128__rotation_3.finished) #(1);
  start__rotator_left_tc__width_128__rotation_4 = 1;
  while(!rotator_left_tc__width_128__rotation_4.finished) #(1);
  start__rotator_left_tc__width_128__rotation_5 = 1;
  while(!rotator_left_tc__width_128__rotation_5.finished) #(1);
  start__rotator_left_tc__width_128__rotation_6 = 1;
  while(!rotator_left_tc__width_128__rotation_6.finished) #(1);
  start__rotator_left_tc__width_128__rotation_7 = 1;
  while(!rotator_left_tc__width_128__rotation_7.finished) #(1);
  start__rotator_left_tc__width_128__rotation_64 = 1;
  while(!rotator_left_tc__width_128__rotation_64.finished) #(1);
  start__rotator_left_tc__width_128__rotation_127 = 1;
  while(!rotator_left_tc__width_128__rotation_127.finished) #(1);
  start__rotator_left_tc__width_128__rotation_128 = 1;
  while(!rotator_left_tc__width_128__rotation_128.finished) #(1);
  start__rotator_left_tc__width_128__rotation_129 = 1;
  while(!rotator_left_tc__width_128__rotation_129.finished) #(1);
  start__rotator_left_tc__width_128__rotation_192 = 1;
  while(!rotator_left_tc__width_128__rotation_192.finished) #(1);
  start__rotator_left_tc__width_128__rotation_255 = 1;
  while(!rotator_left_tc__width_128__rotation_255.finished) #(1);
  start__rotator_left_tc__width_128__rotation_256 = 1;
  while(!rotator_left_tc__width_128__rotation_256.finished) #(1);

  start__rotator_left_tc__width_256__rotation_0 = 1;
  while(!rotator_left_tc__width_256__rotation_0.finished) #(1);
  start__rotator_left_tc__width_256__rotation_1 = 1;
  while(!rotator_left_tc__width_256__rotation_1.finished) #(1);
  start__rotator_left_tc__width_256__rotation_2 = 1;
  while(!rotator_left_tc__width_256__rotation_2.finished) #(1);
  start__rotator_left_tc__width_256__rotation_3 = 1;
  while(!rotator_left_tc__width_256__rotation_3.finished) #(1);
  start__rotator_left_tc__width_256__rotation_4 = 1;
  while(!rotator_left_tc__width_256__rotation_4.finished) #(1);
  start__rotator_left_tc__width_256__rotation_5 = 1;
  while(!rotator_left_tc__width_256__rotation_5.finished) #(1);
  start__rotator_left_tc__width_256__rotation_6 = 1;
  while(!rotator_left_tc__width_256__rotation_6.finished) #(1);
  start__rotator_left_tc__width_256__rotation_7 = 1;
  while(!rotator_left_tc__width_256__rotation_7.finished) #(1);
  start__rotator_left_tc__width_256__rotation_128 = 1;
  while(!rotator_left_tc__width_256__rotation_128.finished) #(1);
  start__rotator_left_tc__width_256__rotation_255 = 1;
  while(!rotator_left_tc__width_256__rotation_255.finished) #(1);
  start__rotator_left_tc__width_256__rotation_256 = 1;
  while(!rotator_left_tc__width_256__rotation_256.finished) #(1);
  start__rotator_left_tc__width_256__rotation_257 = 1;
  while(!rotator_left_tc__width_256__rotation_257.finished) #(1);
  start__rotator_left_tc__width_256__rotation_384 = 1;
  while(!rotator_left_tc__width_256__rotation_384.finished) #(1);
  start__rotator_left_tc__width_256__rotation_511 = 1;
  while(!rotator_left_tc__width_256__rotation_511.finished) #(1);
  start__rotator_left_tc__width_256__rotation_512 = 1;
  while(!rotator_left_tc__width_256__rotation_512.finished) #(1);

  start__rotator_left_tc__width_512__rotation_0 = 1;
  while(!rotator_left_tc__width_512__rotation_0.finished) #(1);
  start__rotator_left_tc__width_512__rotation_1 = 1;
  while(!rotator_left_tc__width_512__rotation_1.finished) #(1);
  start__rotator_left_tc__width_512__rotation_2 = 1;
  while(!rotator_left_tc__width_512__rotation_2.finished) #(1);
  start__rotator_left_tc__width_512__rotation_3 = 1;
  while(!rotator_left_tc__width_512__rotation_3.finished) #(1);
  start__rotator_left_tc__width_512__rotation_4 = 1;
  while(!rotator_left_tc__width_512__rotation_4.finished) #(1);
  start__rotator_left_tc__width_512__rotation_5 = 1;
  while(!rotator_left_tc__width_512__rotation_5.finished) #(1);
  start__rotator_left_tc__width_512__rotation_6 = 1;
  while(!rotator_left_tc__width_512__rotation_6.finished) #(1);
  start__rotator_left_tc__width_512__rotation_7 = 1;
  while(!rotator_left_tc__width_512__rotation_7.finished) #(1);
  start__rotator_left_tc__width_512__rotation_256 = 1;
  while(!rotator_left_tc__width_512__rotation_256.finished) #(1);
  start__rotator_left_tc__width_512__rotation_511 = 1;
  while(!rotator_left_tc__width_512__rotation_511.finished) #(1);
  start__rotator_left_tc__width_512__rotation_512 = 1;
  while(!rotator_left_tc__width_512__rotation_512.finished) #(1);
  start__rotator_left_tc__width_512__rotation_513 = 1;
  while(!rotator_left_tc__width_512__rotation_513.finished) #(1);
  start__rotator_left_tc__width_512__rotation_768 = 1;
  while(!rotator_left_tc__width_512__rotation_768.finished) #(1);
  start__rotator_left_tc__width_512__rotation_1023 = 1;
  while(!rotator_left_tc__width_512__rotation_1023.finished) #(1);
  start__rotator_left_tc__width_512__rotation_1024 = 1;
  while(!rotator_left_tc__width_512__rotation_1024.finished) #(1);

  start__rotator_left_tc__width_1024__rotation_0 = 1;
  while(!rotator_left_tc__width_1024__rotation_0.finished) #(1);
  start__rotator_left_tc__width_1024__rotation_1 = 1;
  while(!rotator_left_tc__width_1024__rotation_1.finished) #(1);
  start__rotator_left_tc__width_1024__rotation_2 = 1;
  while(!rotator_left_tc__width_1024__rotation_2.finished) #(1);
  start__rotator_left_tc__width_1024__rotation_3 = 1;
  while(!rotator_left_tc__width_1024__rotation_3.finished) #(1);
  start__rotator_left_tc__width_1024__rotation_4 = 1;
  while(!rotator_left_tc__width_1024__rotation_4.finished) #(1);
  start__rotator_left_tc__width_1024__rotation_5 = 1;
  while(!rotator_left_tc__width_1024__rotation_5.finished) #(1);
  start__rotator_left_tc__width_1024__rotation_6 = 1;
  while(!rotator_left_tc__width_1024__rotation_6.finished) #(1);
  start__rotator_left_tc__width_1024__rotation_7 = 1;
  while(!rotator_left_tc__width_1024__rotation_7.finished) #(1);
  start__rotator_left_tc__width_1024__rotation_512 = 1;
  while(!rotator_left_tc__width_1024__rotation_512.finished) #(1);
  start__rotator_left_tc__width_1024__rotation_1023 = 1;
  while(!rotator_left_tc__width_1024__rotation_1023.finished) #(1);
  start__rotator_left_tc__width_1024__rotation_1024 = 1;
  while(!rotator_left_tc__width_1024__rotation_1024.finished) #(1);
  start__rotator_left_tc__width_1024__rotation_1025 = 1;
  while(!rotator_left_tc__width_1024__rotation_1025.finished) #(1);
  start__rotator_left_tc__width_1024__rotation_1536 = 1;
  while(!rotator_left_tc__width_1024__rotation_1536.finished) #(1);
  start__rotator_left_tc__width_1024__rotation_2047 = 1;
  while(!rotator_left_tc__width_1024__rotation_2047.finished) #(1);
  start__rotator_left_tc__width_1024__rotation_2048 = 1;
  while(!rotator_left_tc__width_1024__rotation_2048.finished) #(1);


  // Finish
  $finish();
end

endmodule